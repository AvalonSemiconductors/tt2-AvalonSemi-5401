magic
tech sky130A
magscale 1 2
timestamp 1667177658
<< viali >>
rect 1501 20553 1535 20587
rect 1685 20417 1719 20451
rect 1501 18921 1535 18955
rect 2145 18921 2179 18955
rect 1685 18717 1719 18751
rect 2329 18717 2363 18751
rect 1685 18241 1719 18275
rect 2329 18241 2363 18275
rect 1501 18037 1535 18071
rect 2145 18037 2179 18071
rect 2329 17833 2363 17867
rect 2973 17833 3007 17867
rect 1409 17629 1443 17663
rect 2145 17629 2179 17663
rect 3157 17629 3191 17663
rect 1593 17493 1627 17527
rect 2513 17289 2547 17323
rect 3709 17289 3743 17323
rect 2145 17153 2179 17187
rect 3249 17153 3283 17187
rect 3893 17153 3927 17187
rect 1961 17085 1995 17119
rect 2053 17085 2087 17119
rect 3065 16949 3099 16983
rect 1869 16609 1903 16643
rect 3249 16609 3283 16643
rect 4077 16541 4111 16575
rect 4721 16541 4755 16575
rect 2881 16473 2915 16507
rect 3065 16473 3099 16507
rect 1961 16405 1995 16439
rect 2053 16405 2087 16439
rect 2421 16405 2455 16439
rect 3893 16405 3927 16439
rect 4537 16405 4571 16439
rect 4537 16201 4571 16235
rect 2522 16065 2556 16099
rect 4721 16065 4755 16099
rect 5825 16065 5859 16099
rect 2789 15997 2823 16031
rect 3801 15997 3835 16031
rect 4077 15997 4111 16031
rect 4813 15997 4847 16031
rect 5181 15997 5215 16031
rect 1409 15861 1443 15895
rect 5641 15861 5675 15895
rect 5089 15657 5123 15691
rect 3157 15589 3191 15623
rect 5365 15521 5399 15555
rect 5457 15521 5491 15555
rect 1777 15453 1811 15487
rect 4353 15453 4387 15487
rect 4629 15453 4663 15487
rect 5273 15453 5307 15487
rect 5549 15453 5583 15487
rect 6285 15453 6319 15487
rect 2044 15385 2078 15419
rect 6101 15317 6135 15351
rect 5641 15113 5675 15147
rect 3884 15045 3918 15079
rect 6561 15045 6595 15079
rect 2044 14977 2078 15011
rect 5733 14977 5767 15011
rect 5825 14977 5859 15011
rect 6377 14977 6411 15011
rect 6653 14977 6687 15011
rect 7113 14977 7147 15011
rect 1777 14909 1811 14943
rect 3617 14909 3651 14943
rect 5457 14909 5491 14943
rect 6377 14841 6411 14875
rect 3157 14773 3191 14807
rect 4997 14773 5031 14807
rect 5549 14773 5583 14807
rect 7297 14773 7331 14807
rect 2789 14569 2823 14603
rect 6837 14569 6871 14603
rect 5641 14501 5675 14535
rect 7941 14501 7975 14535
rect 6101 14433 6135 14467
rect 6285 14433 6319 14467
rect 1409 14365 1443 14399
rect 5181 14365 5215 14399
rect 7021 14365 7055 14399
rect 7297 14365 7331 14399
rect 7481 14365 7515 14399
rect 8125 14365 8159 14399
rect 1676 14297 1710 14331
rect 4914 14297 4948 14331
rect 3801 14229 3835 14263
rect 6009 14229 6043 14263
rect 3157 14025 3191 14059
rect 6745 14025 6779 14059
rect 8493 14025 8527 14059
rect 1777 13889 1811 13923
rect 2044 13889 2078 13923
rect 3617 13889 3651 13923
rect 3884 13889 3918 13923
rect 5549 13889 5583 13923
rect 5641 13889 5675 13923
rect 7629 13889 7663 13923
rect 7757 13889 7791 13923
rect 7849 13889 7883 13923
rect 8677 13889 8711 13923
rect 9321 13889 9355 13923
rect 6837 13821 6871 13855
rect 6929 13821 6963 13855
rect 8033 13821 8067 13855
rect 4997 13753 5031 13787
rect 5825 13753 5859 13787
rect 6377 13753 6411 13787
rect 9137 13685 9171 13719
rect 3065 13481 3099 13515
rect 5181 13481 5215 13515
rect 9689 13413 9723 13447
rect 7941 13345 7975 13379
rect 8033 13345 8067 13379
rect 9045 13345 9079 13379
rect 1685 13277 1719 13311
rect 3801 13277 3835 13311
rect 7021 13277 7055 13311
rect 7849 13277 7883 13311
rect 8953 13277 8987 13311
rect 9873 13277 9907 13311
rect 1930 13209 1964 13243
rect 4068 13209 4102 13243
rect 6754 13209 6788 13243
rect 9229 13209 9263 13243
rect 5641 13141 5675 13175
rect 7481 13141 7515 13175
rect 8953 13141 8987 13175
rect 1409 12937 1443 12971
rect 5733 12937 5767 12971
rect 8677 12869 8711 12903
rect 9321 12869 9355 12903
rect 1593 12801 1627 12835
rect 2697 12801 2731 12835
rect 2973 12801 3007 12835
rect 3893 12801 3927 12835
rect 4353 12801 4387 12835
rect 4620 12801 4654 12835
rect 7490 12801 7524 12835
rect 7757 12801 7791 12835
rect 8401 12801 8435 12835
rect 9505 12801 9539 12835
rect 9965 12801 9999 12835
rect 10609 12801 10643 12835
rect 2053 12733 2087 12767
rect 2856 12733 2890 12767
rect 3709 12733 3743 12767
rect 8585 12733 8619 12767
rect 3249 12665 3283 12699
rect 9137 12665 9171 12699
rect 6377 12597 6411 12631
rect 8217 12597 8251 12631
rect 8401 12597 8435 12631
rect 10057 12597 10091 12631
rect 10793 12597 10827 12631
rect 1409 12393 1443 12427
rect 7941 12393 7975 12427
rect 8309 12393 8343 12427
rect 10793 12393 10827 12427
rect 11345 12393 11379 12427
rect 12081 12393 12115 12427
rect 2605 12325 2639 12359
rect 6101 12325 6135 12359
rect 8953 12325 8987 12359
rect 2191 12257 2225 12291
rect 2329 12257 2363 12291
rect 3249 12257 3283 12291
rect 4445 12257 4479 12291
rect 4604 12257 4638 12291
rect 4997 12257 5031 12291
rect 5457 12257 5491 12291
rect 10701 12257 10735 12291
rect 2053 12189 2087 12223
rect 3065 12189 3099 12223
rect 4721 12189 4755 12223
rect 5641 12189 5675 12223
rect 7481 12189 7515 12223
rect 8125 12189 8159 12223
rect 8217 12189 8251 12223
rect 9137 12189 9171 12223
rect 9229 12189 9263 12223
rect 9321 12189 9355 12223
rect 10057 12189 10091 12223
rect 10609 12189 10643 12223
rect 11529 12189 11563 12223
rect 11989 12189 12023 12223
rect 12173 12189 12207 12223
rect 7236 12121 7270 12155
rect 8401 12121 8435 12155
rect 10885 12121 10919 12155
rect 3801 12053 3835 12087
rect 9965 12053 9999 12087
rect 1869 11849 1903 11883
rect 4169 11849 4203 11883
rect 8217 11849 8251 11883
rect 5282 11781 5316 11815
rect 10333 11781 10367 11815
rect 5549 11713 5583 11747
rect 7490 11713 7524 11747
rect 7757 11713 7791 11747
rect 8585 11713 8619 11747
rect 9505 11713 9539 11747
rect 10517 11713 10551 11747
rect 11713 11713 11747 11747
rect 12173 11713 12207 11747
rect 12357 11713 12391 11747
rect 2513 11645 2547 11679
rect 2672 11645 2706 11679
rect 2789 11645 2823 11679
rect 3525 11645 3559 11679
rect 3709 11645 3743 11679
rect 8677 11645 8711 11679
rect 9597 11645 9631 11679
rect 9689 11645 9723 11679
rect 9781 11645 9815 11679
rect 10793 11645 10827 11679
rect 3065 11577 3099 11611
rect 6377 11509 6411 11543
rect 8861 11509 8895 11543
rect 9321 11509 9355 11543
rect 10701 11509 10735 11543
rect 11529 11509 11563 11543
rect 12265 11509 12299 11543
rect 1455 11305 1489 11339
rect 3801 11305 3835 11339
rect 5641 11305 5675 11339
rect 7481 11305 7515 11339
rect 9689 11305 9723 11339
rect 10149 11305 10183 11339
rect 11621 11305 11655 11339
rect 13369 11237 13403 11271
rect 2881 11169 2915 11203
rect 5181 11169 5215 11203
rect 8033 11169 8067 11203
rect 9045 11169 9079 11203
rect 3249 11101 3283 11135
rect 7021 11101 7055 11135
rect 10333 11101 10367 11135
rect 10701 11101 10735 11135
rect 11161 11101 11195 11135
rect 11437 11101 11471 11135
rect 12265 11101 12299 11135
rect 12909 11101 12943 11135
rect 13553 11101 13587 11135
rect 4936 11033 4970 11067
rect 6776 11033 6810 11067
rect 9321 11033 9355 11067
rect 10425 11033 10459 11067
rect 10517 11033 10551 11067
rect 7849 10965 7883 10999
rect 7941 10965 7975 10999
rect 9229 10965 9263 10999
rect 11253 10965 11287 10999
rect 12081 10965 12115 10999
rect 12725 10965 12759 10999
rect 3617 10761 3651 10795
rect 9597 10761 9631 10795
rect 11529 10761 11563 10795
rect 4730 10693 4764 10727
rect 5457 10693 5491 10727
rect 5673 10693 5707 10727
rect 8484 10693 8518 10727
rect 13921 10693 13955 10727
rect 6633 10625 6667 10659
rect 8217 10625 8251 10659
rect 10333 10625 10367 10659
rect 10425 10625 10459 10659
rect 11713 10625 11747 10659
rect 12449 10625 12483 10659
rect 12541 10625 12575 10659
rect 12725 10625 12759 10659
rect 13185 10625 13219 10659
rect 13369 10625 13403 10659
rect 13829 10625 13863 10659
rect 14013 10625 14047 10659
rect 14657 10625 14691 10659
rect 1409 10557 1443 10591
rect 1685 10557 1719 10591
rect 4997 10557 5031 10591
rect 6377 10557 6411 10591
rect 10241 10557 10275 10591
rect 10517 10557 10551 10591
rect 11989 10557 12023 10591
rect 7757 10489 7791 10523
rect 11897 10489 11931 10523
rect 13185 10489 13219 10523
rect 3157 10421 3191 10455
rect 5641 10421 5675 10455
rect 5825 10421 5859 10455
rect 10057 10421 10091 10455
rect 12725 10421 12759 10455
rect 14473 10421 14507 10455
rect 3801 10217 3835 10251
rect 8125 10217 8159 10251
rect 10793 10217 10827 10251
rect 14105 10217 14139 10251
rect 7021 10149 7055 10183
rect 11253 10149 11287 10183
rect 13185 10149 13219 10183
rect 5181 10081 5215 10115
rect 5641 10081 5675 10115
rect 9045 10081 9079 10115
rect 11529 10081 11563 10115
rect 1501 10013 1535 10047
rect 4914 10013 4948 10047
rect 7481 10013 7515 10047
rect 7629 10013 7663 10047
rect 7757 10013 7791 10047
rect 7987 10013 8021 10047
rect 10149 10013 10183 10047
rect 10333 10013 10367 10047
rect 10425 10013 10459 10047
rect 10563 10013 10597 10047
rect 11621 10013 11655 10047
rect 12265 10013 12299 10047
rect 12357 10013 12391 10047
rect 12541 10013 12575 10047
rect 13369 10013 13403 10047
rect 14289 10013 14323 10047
rect 1777 9945 1811 9979
rect 5886 9945 5920 9979
rect 7849 9945 7883 9979
rect 9321 9945 9355 9979
rect 3249 9877 3283 9911
rect 9229 9877 9263 9911
rect 9689 9877 9723 9911
rect 12725 9877 12759 9911
rect 1593 9673 1627 9707
rect 13277 9673 13311 9707
rect 5273 9605 5307 9639
rect 9873 9605 9907 9639
rect 10609 9605 10643 9639
rect 6644 9537 6678 9571
rect 8493 9537 8527 9571
rect 8861 9537 8895 9571
rect 9505 9537 9539 9571
rect 9597 9517 9631 9551
rect 10425 9537 10459 9571
rect 10701 9537 10735 9571
rect 10793 9537 10827 9571
rect 11713 9537 11747 9571
rect 12357 9537 12391 9571
rect 12541 9537 12575 9571
rect 12633 9537 12667 9571
rect 13093 9537 13127 9571
rect 13277 9537 13311 9571
rect 3065 9469 3099 9503
rect 3341 9469 3375 9503
rect 5549 9469 5583 9503
rect 6377 9469 6411 9503
rect 8401 9469 8435 9503
rect 9965 9469 9999 9503
rect 11529 9469 11563 9503
rect 11897 9469 11931 9503
rect 7757 9401 7791 9435
rect 8217 9401 8251 9435
rect 10977 9401 11011 9435
rect 12449 9401 12483 9435
rect 3801 9333 3835 9367
rect 9321 9333 9355 9367
rect 1455 9129 1489 9163
rect 7849 9129 7883 9163
rect 10149 9129 10183 9163
rect 12541 9129 12575 9163
rect 5549 9061 5583 9095
rect 7757 9061 7791 9095
rect 3801 8993 3835 9027
rect 6285 8993 6319 9027
rect 11161 8993 11195 9027
rect 2881 8925 2915 8959
rect 3249 8925 3283 8959
rect 6009 8925 6043 8959
rect 7573 8925 7607 8959
rect 7665 8925 7699 8959
rect 8033 8925 8067 8959
rect 9137 8925 9171 8959
rect 9321 8925 9355 8959
rect 9505 8925 9539 8959
rect 10517 8925 10551 8959
rect 10977 8925 11011 8959
rect 11345 8925 11379 8959
rect 11989 8925 12023 8959
rect 12449 8925 12483 8959
rect 12633 8925 12667 8959
rect 4077 8857 4111 8891
rect 9229 8857 9263 8891
rect 7297 8789 7331 8823
rect 8953 8789 8987 8823
rect 9965 8789 9999 8823
rect 10149 8789 10183 8823
rect 11069 8789 11103 8823
rect 11253 8789 11287 8823
rect 11805 8789 11839 8823
rect 7113 8585 7147 8619
rect 9781 8585 9815 8619
rect 11713 8585 11747 8619
rect 12173 8585 12207 8619
rect 3203 8517 3237 8551
rect 3985 8517 4019 8551
rect 8217 8517 8251 8551
rect 3709 8449 3743 8483
rect 6653 8449 6687 8483
rect 6745 8449 6779 8483
rect 7849 8449 7883 8483
rect 8125 8449 8159 8483
rect 8953 8449 8987 8483
rect 9229 8449 9263 8483
rect 9689 8449 9723 8483
rect 9945 8449 9979 8483
rect 10609 8449 10643 8483
rect 10793 8449 10827 8483
rect 11529 8449 11563 8483
rect 12173 8449 12207 8483
rect 12357 8449 12391 8483
rect 1409 8381 1443 8415
rect 1777 8381 1811 8415
rect 6561 8381 6595 8415
rect 7757 8381 7791 8415
rect 10977 8381 11011 8415
rect 5457 8313 5491 8347
rect 7573 8313 7607 8347
rect 8677 8313 8711 8347
rect 10149 8313 10183 8347
rect 9137 8245 9171 8279
rect 3157 8041 3191 8075
rect 5549 8041 5583 8075
rect 7573 8041 7607 8075
rect 7757 8041 7791 8075
rect 8309 8041 8343 8075
rect 10057 8041 10091 8075
rect 11897 8041 11931 8075
rect 6745 7973 6779 8007
rect 9045 7973 9079 8007
rect 6193 7905 6227 7939
rect 11253 7905 11287 7939
rect 1409 7837 1443 7871
rect 3801 7837 3835 7871
rect 7205 7837 7239 7871
rect 8401 7837 8435 7871
rect 9873 7837 9907 7871
rect 10517 7837 10551 7871
rect 10701 7837 10735 7871
rect 11161 7837 11195 7871
rect 11345 7837 11379 7871
rect 11805 7837 11839 7871
rect 11989 7837 12023 7871
rect 1685 7769 1719 7803
rect 4077 7769 4111 7803
rect 9413 7769 9447 7803
rect 6285 7701 6319 7735
rect 6377 7701 6411 7735
rect 7573 7701 7607 7735
rect 8953 7701 8987 7735
rect 10609 7701 10643 7735
rect 6929 7497 6963 7531
rect 8769 7497 8803 7531
rect 10517 7497 10551 7531
rect 6653 7429 6687 7463
rect 8401 7429 8435 7463
rect 1501 7361 1535 7395
rect 3976 7361 4010 7395
rect 5549 7361 5583 7395
rect 5641 7361 5675 7395
rect 5828 7361 5862 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 6769 7361 6803 7395
rect 7573 7361 7607 7395
rect 8585 7361 8619 7395
rect 9237 7359 9271 7393
rect 9423 7361 9457 7395
rect 9873 7361 9907 7395
rect 10057 7361 10091 7395
rect 10517 7361 10551 7395
rect 10701 7361 10735 7395
rect 1777 7293 1811 7327
rect 3709 7293 3743 7327
rect 7481 7293 7515 7327
rect 7941 7293 7975 7327
rect 5089 7225 5123 7259
rect 5825 7225 5859 7259
rect 3249 7157 3283 7191
rect 9321 7157 9355 7191
rect 9965 7157 9999 7191
rect 1666 6953 1700 6987
rect 3157 6953 3191 6987
rect 5181 6953 5215 6987
rect 5641 6953 5675 6987
rect 6101 6953 6135 6987
rect 9045 6953 9079 6987
rect 9597 6953 9631 6987
rect 1409 6817 1443 6851
rect 3801 6817 3835 6851
rect 4077 6817 4111 6851
rect 5365 6817 5399 6851
rect 6285 6817 6319 6851
rect 7573 6817 7607 6851
rect 5089 6749 5123 6783
rect 6101 6749 6135 6783
rect 6377 6749 6411 6783
rect 7113 6749 7147 6783
rect 7205 6749 7239 6783
rect 7389 6749 7423 6783
rect 8033 6749 8067 6783
rect 8217 6749 8251 6783
rect 8309 6749 8343 6783
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 9597 6749 9631 6783
rect 9781 6749 9815 6783
rect 6561 6613 6595 6647
rect 2789 6409 2823 6443
rect 5089 6409 5123 6443
rect 5733 6409 5767 6443
rect 6377 6409 6411 6443
rect 7297 6409 7331 6443
rect 8309 6409 8343 6443
rect 1676 6341 1710 6375
rect 4721 6341 4755 6375
rect 4813 6341 4847 6375
rect 5549 6341 5583 6375
rect 7449 6341 7483 6375
rect 7665 6341 7699 6375
rect 1409 6273 1443 6307
rect 3801 6273 3835 6307
rect 4537 6273 4571 6307
rect 4905 6273 4939 6307
rect 5809 6273 5843 6307
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 6837 6273 6871 6307
rect 8125 6273 8159 6307
rect 8953 6273 8987 6307
rect 4077 6205 4111 6239
rect 5549 6137 5583 6171
rect 8769 6137 8803 6171
rect 7490 6069 7524 6103
rect 6285 5865 6319 5899
rect 7665 5865 7699 5899
rect 4077 5729 4111 5763
rect 5181 5729 5215 5763
rect 5641 5729 5675 5763
rect 7021 5729 7055 5763
rect 2421 5661 2455 5695
rect 2697 5661 2731 5695
rect 3801 5661 3835 5695
rect 5273 5661 5307 5695
rect 6929 5661 6963 5695
rect 7113 5661 7147 5695
rect 7573 5661 7607 5695
rect 7757 5661 7791 5695
rect 8401 5661 8435 5695
rect 6101 5593 6135 5627
rect 6301 5525 6335 5559
rect 6469 5525 6503 5559
rect 8217 5525 8251 5559
rect 3617 5321 3651 5355
rect 5089 5321 5123 5355
rect 6469 5321 6503 5355
rect 3341 5253 3375 5287
rect 5457 5253 5491 5287
rect 5227 5219 5261 5253
rect 2329 5185 2363 5219
rect 3065 5185 3099 5219
rect 3249 5185 3283 5219
rect 3433 5185 3467 5219
rect 4261 5185 4295 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 7021 5185 7055 5219
rect 2605 5117 2639 5151
rect 4353 5117 4387 5151
rect 7205 5049 7239 5083
rect 4629 4981 4663 5015
rect 5273 4981 5307 5015
rect 3065 4777 3099 4811
rect 4261 4777 4295 4811
rect 6101 4777 6135 4811
rect 6837 4777 6871 4811
rect 2697 4709 2731 4743
rect 3249 4709 3283 4743
rect 1409 4641 1443 4675
rect 1685 4641 1719 4675
rect 5457 4641 5491 4675
rect 3801 4573 3835 4607
rect 4077 4573 4111 4607
rect 4721 4573 4755 4607
rect 5365 4573 5399 4607
rect 6009 4573 6043 4607
rect 6193 4573 6227 4607
rect 6653 4573 6687 4607
rect 3893 4505 3927 4539
rect 3065 4437 3099 4471
rect 4905 4437 4939 4471
rect 2697 4233 2731 4267
rect 3617 4165 3651 4199
rect 3801 4165 3835 4199
rect 1685 4097 1719 4131
rect 2881 4097 2915 4131
rect 3065 4097 3099 4131
rect 3157 4097 3191 4131
rect 4629 4097 4663 4131
rect 5089 4097 5123 4131
rect 5273 4097 5307 4131
rect 1409 4029 1443 4063
rect 3985 4029 4019 4063
rect 5181 3961 5215 3995
rect 4537 3893 4571 3927
rect 3893 3689 3927 3723
rect 3065 3621 3099 3655
rect 4445 3621 4479 3655
rect 2329 3553 2363 3587
rect 1501 3485 1535 3519
rect 1685 3485 1719 3519
rect 2145 3485 2179 3519
rect 2237 3485 2271 3519
rect 2513 3485 2547 3519
rect 2973 3485 3007 3519
rect 3157 3485 3191 3519
rect 3801 3485 3835 3519
rect 3985 3485 4019 3519
rect 4629 3485 4663 3519
rect 1593 3417 1627 3451
rect 2421 3349 2455 3383
rect 2421 3145 2455 3179
rect 3065 3145 3099 3179
rect 1501 3009 1535 3043
rect 2237 3009 2271 3043
rect 2881 3009 2915 3043
rect 3065 3009 3099 3043
rect 3709 3009 3743 3043
rect 3525 2873 3559 2907
rect 1685 2805 1719 2839
rect 2881 2601 2915 2635
rect 1685 2465 1719 2499
rect 1409 2397 1443 2431
rect 2697 2397 2731 2431
rect 1593 2057 1627 2091
rect 1409 1921 1443 1955
rect 2053 1921 2087 1955
rect 2237 1921 2271 1955
rect 2145 1853 2179 1887
rect 1409 1309 1443 1343
rect 1593 1173 1627 1207
<< metal1 >>
rect 1104 22874 16836 22896
rect 1104 22822 4898 22874
rect 4950 22822 4962 22874
rect 5014 22822 5026 22874
rect 5078 22822 5090 22874
rect 5142 22822 5154 22874
rect 5206 22822 8846 22874
rect 8898 22822 8910 22874
rect 8962 22822 8974 22874
rect 9026 22822 9038 22874
rect 9090 22822 9102 22874
rect 9154 22822 12794 22874
rect 12846 22822 12858 22874
rect 12910 22822 12922 22874
rect 12974 22822 12986 22874
rect 13038 22822 13050 22874
rect 13102 22822 16836 22874
rect 1104 22800 16836 22822
rect 1104 22330 16836 22352
rect 1104 22278 2924 22330
rect 2976 22278 2988 22330
rect 3040 22278 3052 22330
rect 3104 22278 3116 22330
rect 3168 22278 3180 22330
rect 3232 22278 6872 22330
rect 6924 22278 6936 22330
rect 6988 22278 7000 22330
rect 7052 22278 7064 22330
rect 7116 22278 7128 22330
rect 7180 22278 10820 22330
rect 10872 22278 10884 22330
rect 10936 22278 10948 22330
rect 11000 22278 11012 22330
rect 11064 22278 11076 22330
rect 11128 22278 14768 22330
rect 14820 22278 14832 22330
rect 14884 22278 14896 22330
rect 14948 22278 14960 22330
rect 15012 22278 15024 22330
rect 15076 22278 16836 22330
rect 1104 22256 16836 22278
rect 1104 21786 16836 21808
rect 1104 21734 4898 21786
rect 4950 21734 4962 21786
rect 5014 21734 5026 21786
rect 5078 21734 5090 21786
rect 5142 21734 5154 21786
rect 5206 21734 8846 21786
rect 8898 21734 8910 21786
rect 8962 21734 8974 21786
rect 9026 21734 9038 21786
rect 9090 21734 9102 21786
rect 9154 21734 12794 21786
rect 12846 21734 12858 21786
rect 12910 21734 12922 21786
rect 12974 21734 12986 21786
rect 13038 21734 13050 21786
rect 13102 21734 16836 21786
rect 1104 21712 16836 21734
rect 1104 21242 16836 21264
rect 1104 21190 2924 21242
rect 2976 21190 2988 21242
rect 3040 21190 3052 21242
rect 3104 21190 3116 21242
rect 3168 21190 3180 21242
rect 3232 21190 6872 21242
rect 6924 21190 6936 21242
rect 6988 21190 7000 21242
rect 7052 21190 7064 21242
rect 7116 21190 7128 21242
rect 7180 21190 10820 21242
rect 10872 21190 10884 21242
rect 10936 21190 10948 21242
rect 11000 21190 11012 21242
rect 11064 21190 11076 21242
rect 11128 21190 14768 21242
rect 14820 21190 14832 21242
rect 14884 21190 14896 21242
rect 14948 21190 14960 21242
rect 15012 21190 15024 21242
rect 15076 21190 16836 21242
rect 1104 21168 16836 21190
rect 1104 20698 16836 20720
rect 1104 20646 4898 20698
rect 4950 20646 4962 20698
rect 5014 20646 5026 20698
rect 5078 20646 5090 20698
rect 5142 20646 5154 20698
rect 5206 20646 8846 20698
rect 8898 20646 8910 20698
rect 8962 20646 8974 20698
rect 9026 20646 9038 20698
rect 9090 20646 9102 20698
rect 9154 20646 12794 20698
rect 12846 20646 12858 20698
rect 12910 20646 12922 20698
rect 12974 20646 12986 20698
rect 13038 20646 13050 20698
rect 13102 20646 16836 20698
rect 1104 20624 16836 20646
rect 1489 20587 1547 20593
rect 1489 20553 1501 20587
rect 1535 20584 1547 20587
rect 2774 20584 2780 20596
rect 1535 20556 2780 20584
rect 1535 20553 1547 20556
rect 1489 20547 1547 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 1670 20448 1676 20460
rect 1631 20420 1676 20448
rect 1670 20408 1676 20420
rect 1728 20408 1734 20460
rect 1104 20154 16836 20176
rect 1104 20102 2924 20154
rect 2976 20102 2988 20154
rect 3040 20102 3052 20154
rect 3104 20102 3116 20154
rect 3168 20102 3180 20154
rect 3232 20102 6872 20154
rect 6924 20102 6936 20154
rect 6988 20102 7000 20154
rect 7052 20102 7064 20154
rect 7116 20102 7128 20154
rect 7180 20102 10820 20154
rect 10872 20102 10884 20154
rect 10936 20102 10948 20154
rect 11000 20102 11012 20154
rect 11064 20102 11076 20154
rect 11128 20102 14768 20154
rect 14820 20102 14832 20154
rect 14884 20102 14896 20154
rect 14948 20102 14960 20154
rect 15012 20102 15024 20154
rect 15076 20102 16836 20154
rect 1104 20080 16836 20102
rect 1104 19610 16836 19632
rect 1104 19558 4898 19610
rect 4950 19558 4962 19610
rect 5014 19558 5026 19610
rect 5078 19558 5090 19610
rect 5142 19558 5154 19610
rect 5206 19558 8846 19610
rect 8898 19558 8910 19610
rect 8962 19558 8974 19610
rect 9026 19558 9038 19610
rect 9090 19558 9102 19610
rect 9154 19558 12794 19610
rect 12846 19558 12858 19610
rect 12910 19558 12922 19610
rect 12974 19558 12986 19610
rect 13038 19558 13050 19610
rect 13102 19558 16836 19610
rect 1104 19536 16836 19558
rect 1104 19066 16836 19088
rect 1104 19014 2924 19066
rect 2976 19014 2988 19066
rect 3040 19014 3052 19066
rect 3104 19014 3116 19066
rect 3168 19014 3180 19066
rect 3232 19014 6872 19066
rect 6924 19014 6936 19066
rect 6988 19014 7000 19066
rect 7052 19014 7064 19066
rect 7116 19014 7128 19066
rect 7180 19014 10820 19066
rect 10872 19014 10884 19066
rect 10936 19014 10948 19066
rect 11000 19014 11012 19066
rect 11064 19014 11076 19066
rect 11128 19014 14768 19066
rect 14820 19014 14832 19066
rect 14884 19014 14896 19066
rect 14948 19014 14960 19066
rect 15012 19014 15024 19066
rect 15076 19014 16836 19066
rect 1104 18992 16836 19014
rect 1486 18952 1492 18964
rect 1447 18924 1492 18952
rect 1486 18912 1492 18924
rect 1544 18912 1550 18964
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 2133 18955 2191 18961
rect 2133 18952 2145 18955
rect 1728 18924 2145 18952
rect 1728 18912 1734 18924
rect 2133 18921 2145 18924
rect 2179 18921 2191 18955
rect 2133 18915 2191 18921
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18717 1731 18751
rect 2314 18748 2320 18760
rect 2275 18720 2320 18748
rect 1673 18711 1731 18717
rect 1688 18680 1716 18711
rect 2314 18708 2320 18720
rect 2372 18708 2378 18760
rect 4798 18680 4804 18692
rect 1688 18652 4804 18680
rect 4798 18640 4804 18652
rect 4856 18640 4862 18692
rect 1104 18522 16836 18544
rect 1104 18470 4898 18522
rect 4950 18470 4962 18522
rect 5014 18470 5026 18522
rect 5078 18470 5090 18522
rect 5142 18470 5154 18522
rect 5206 18470 8846 18522
rect 8898 18470 8910 18522
rect 8962 18470 8974 18522
rect 9026 18470 9038 18522
rect 9090 18470 9102 18522
rect 9154 18470 12794 18522
rect 12846 18470 12858 18522
rect 12910 18470 12922 18522
rect 12974 18470 12986 18522
rect 13038 18470 13050 18522
rect 13102 18470 16836 18522
rect 1104 18448 16836 18470
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 1673 18235 1731 18241
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 2406 18272 2412 18284
rect 2363 18244 2412 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 1688 18204 1716 18235
rect 2406 18232 2412 18244
rect 2464 18232 2470 18284
rect 3694 18204 3700 18216
rect 1688 18176 3700 18204
rect 3694 18164 3700 18176
rect 3752 18164 3758 18216
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 2130 18068 2136 18080
rect 2091 18040 2136 18068
rect 2130 18028 2136 18040
rect 2188 18028 2194 18080
rect 1104 17978 16836 18000
rect 1104 17926 2924 17978
rect 2976 17926 2988 17978
rect 3040 17926 3052 17978
rect 3104 17926 3116 17978
rect 3168 17926 3180 17978
rect 3232 17926 6872 17978
rect 6924 17926 6936 17978
rect 6988 17926 7000 17978
rect 7052 17926 7064 17978
rect 7116 17926 7128 17978
rect 7180 17926 10820 17978
rect 10872 17926 10884 17978
rect 10936 17926 10948 17978
rect 11000 17926 11012 17978
rect 11064 17926 11076 17978
rect 11128 17926 14768 17978
rect 14820 17926 14832 17978
rect 14884 17926 14896 17978
rect 14948 17926 14960 17978
rect 15012 17926 15024 17978
rect 15076 17926 16836 17978
rect 1104 17904 16836 17926
rect 2317 17867 2375 17873
rect 2317 17833 2329 17867
rect 2363 17864 2375 17867
rect 2774 17864 2780 17876
rect 2363 17836 2780 17864
rect 2363 17833 2375 17836
rect 2317 17827 2375 17833
rect 2774 17824 2780 17836
rect 2832 17824 2838 17876
rect 2961 17867 3019 17873
rect 2961 17833 2973 17867
rect 3007 17864 3019 17867
rect 3326 17864 3332 17876
rect 3007 17836 3332 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 3326 17824 3332 17836
rect 3384 17824 3390 17876
rect 1394 17660 1400 17672
rect 1355 17632 1400 17660
rect 1394 17620 1400 17632
rect 1452 17620 1458 17672
rect 2130 17660 2136 17672
rect 2091 17632 2136 17660
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 3145 17663 3203 17669
rect 3145 17629 3157 17663
rect 3191 17660 3203 17663
rect 4522 17660 4528 17672
rect 3191 17632 4528 17660
rect 3191 17629 3203 17632
rect 3145 17623 3203 17629
rect 4522 17620 4528 17632
rect 4580 17620 4586 17672
rect 3326 17592 3332 17604
rect 1596 17564 3332 17592
rect 1596 17533 1624 17564
rect 3326 17552 3332 17564
rect 3384 17552 3390 17604
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17493 1639 17527
rect 1581 17487 1639 17493
rect 1104 17434 16836 17456
rect 1104 17382 4898 17434
rect 4950 17382 4962 17434
rect 5014 17382 5026 17434
rect 5078 17382 5090 17434
rect 5142 17382 5154 17434
rect 5206 17382 8846 17434
rect 8898 17382 8910 17434
rect 8962 17382 8974 17434
rect 9026 17382 9038 17434
rect 9090 17382 9102 17434
rect 9154 17382 12794 17434
rect 12846 17382 12858 17434
rect 12910 17382 12922 17434
rect 12974 17382 12986 17434
rect 13038 17382 13050 17434
rect 13102 17382 16836 17434
rect 1104 17360 16836 17382
rect 2314 17280 2320 17332
rect 2372 17320 2378 17332
rect 2501 17323 2559 17329
rect 2501 17320 2513 17323
rect 2372 17292 2513 17320
rect 2372 17280 2378 17292
rect 2501 17289 2513 17292
rect 2547 17289 2559 17323
rect 3694 17320 3700 17332
rect 3655 17292 3700 17320
rect 2501 17283 2559 17289
rect 3694 17280 3700 17292
rect 3752 17280 3758 17332
rect 11330 17252 11336 17264
rect 3252 17224 11336 17252
rect 3252 17193 3280 17224
rect 11330 17212 11336 17224
rect 11388 17212 11394 17264
rect 2133 17187 2191 17193
rect 2133 17184 2145 17187
rect 1504 17156 2145 17184
rect 1504 17128 1532 17156
rect 2133 17153 2145 17156
rect 2179 17153 2191 17187
rect 2133 17147 2191 17153
rect 3237 17187 3295 17193
rect 3237 17153 3249 17187
rect 3283 17153 3295 17187
rect 3237 17147 3295 17153
rect 3881 17187 3939 17193
rect 3881 17153 3893 17187
rect 3927 17153 3939 17187
rect 3881 17147 3939 17153
rect 1486 17076 1492 17128
rect 1544 17076 1550 17128
rect 1946 17116 1952 17128
rect 1907 17088 1952 17116
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 2056 17048 2084 17079
rect 2314 17076 2320 17128
rect 2372 17116 2378 17128
rect 3896 17116 3924 17147
rect 2372 17088 3924 17116
rect 2372 17076 2378 17088
rect 6270 17048 6276 17060
rect 2056 17020 6276 17048
rect 6270 17008 6276 17020
rect 6328 17008 6334 17060
rect 3053 16983 3111 16989
rect 3053 16949 3065 16983
rect 3099 16980 3111 16983
rect 3510 16980 3516 16992
rect 3099 16952 3516 16980
rect 3099 16949 3111 16952
rect 3053 16943 3111 16949
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 1104 16890 16836 16912
rect 1104 16838 2924 16890
rect 2976 16838 2988 16890
rect 3040 16838 3052 16890
rect 3104 16838 3116 16890
rect 3168 16838 3180 16890
rect 3232 16838 6872 16890
rect 6924 16838 6936 16890
rect 6988 16838 7000 16890
rect 7052 16838 7064 16890
rect 7116 16838 7128 16890
rect 7180 16838 10820 16890
rect 10872 16838 10884 16890
rect 10936 16838 10948 16890
rect 11000 16838 11012 16890
rect 11064 16838 11076 16890
rect 11128 16838 14768 16890
rect 14820 16838 14832 16890
rect 14884 16838 14896 16890
rect 14948 16838 14960 16890
rect 15012 16838 15024 16890
rect 15076 16838 16836 16890
rect 1104 16816 16836 16838
rect 1946 16708 1952 16720
rect 1859 16680 1952 16708
rect 1872 16649 1900 16680
rect 1946 16668 1952 16680
rect 2004 16708 2010 16720
rect 4338 16708 4344 16720
rect 2004 16680 4344 16708
rect 2004 16668 2010 16680
rect 4338 16668 4344 16680
rect 4396 16668 4402 16720
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16609 1915 16643
rect 1857 16603 1915 16609
rect 3237 16643 3295 16649
rect 3237 16609 3249 16643
rect 3283 16640 3295 16643
rect 9214 16640 9220 16652
rect 3283 16612 9220 16640
rect 3283 16609 3295 16612
rect 3237 16603 3295 16609
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 4706 16572 4712 16584
rect 4667 16544 4712 16572
rect 4065 16535 4123 16541
rect 2498 16464 2504 16516
rect 2556 16504 2562 16516
rect 2869 16507 2927 16513
rect 2869 16504 2881 16507
rect 2556 16476 2881 16504
rect 2556 16464 2562 16476
rect 2869 16473 2881 16476
rect 2915 16473 2927 16507
rect 3050 16504 3056 16516
rect 3011 16476 3056 16504
rect 2869 16467 2927 16473
rect 3050 16464 3056 16476
rect 3108 16464 3114 16516
rect 4080 16504 4108 16535
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 6730 16504 6736 16516
rect 3160 16476 3924 16504
rect 4080 16476 6736 16504
rect 1946 16436 1952 16448
rect 1907 16408 1952 16436
rect 1946 16396 1952 16408
rect 2004 16396 2010 16448
rect 2038 16396 2044 16448
rect 2096 16436 2102 16448
rect 2406 16436 2412 16448
rect 2096 16408 2141 16436
rect 2367 16408 2412 16436
rect 2096 16396 2102 16408
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 3160 16436 3188 16476
rect 3896 16445 3924 16476
rect 6730 16464 6736 16476
rect 6788 16464 6794 16516
rect 2832 16408 3188 16436
rect 3881 16439 3939 16445
rect 2832 16396 2838 16408
rect 3881 16405 3893 16439
rect 3927 16405 3939 16439
rect 3881 16399 3939 16405
rect 3970 16396 3976 16448
rect 4028 16436 4034 16448
rect 4525 16439 4583 16445
rect 4525 16436 4537 16439
rect 4028 16408 4537 16436
rect 4028 16396 4034 16408
rect 4525 16405 4537 16408
rect 4571 16405 4583 16439
rect 4525 16399 4583 16405
rect 1104 16346 16836 16368
rect 1104 16294 4898 16346
rect 4950 16294 4962 16346
rect 5014 16294 5026 16346
rect 5078 16294 5090 16346
rect 5142 16294 5154 16346
rect 5206 16294 8846 16346
rect 8898 16294 8910 16346
rect 8962 16294 8974 16346
rect 9026 16294 9038 16346
rect 9090 16294 9102 16346
rect 9154 16294 12794 16346
rect 12846 16294 12858 16346
rect 12910 16294 12922 16346
rect 12974 16294 12986 16346
rect 13038 16294 13050 16346
rect 13102 16294 16836 16346
rect 1104 16272 16836 16294
rect 4522 16232 4528 16244
rect 4483 16204 4528 16232
rect 4522 16192 4528 16204
rect 4580 16192 4586 16244
rect 1670 16056 1676 16108
rect 1728 16096 1734 16108
rect 2510 16099 2568 16105
rect 2510 16096 2522 16099
rect 1728 16068 2522 16096
rect 1728 16056 1734 16068
rect 2510 16065 2522 16068
rect 2556 16065 2568 16099
rect 2510 16059 2568 16065
rect 4709 16099 4767 16105
rect 4709 16065 4721 16099
rect 4755 16096 4767 16099
rect 5442 16096 5448 16108
rect 4755 16068 5448 16096
rect 4755 16065 4767 16068
rect 4709 16059 4767 16065
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 5810 16096 5816 16108
rect 5771 16068 5816 16096
rect 5810 16056 5816 16068
rect 5868 16056 5874 16108
rect 2777 16031 2835 16037
rect 2777 15997 2789 16031
rect 2823 16028 2835 16031
rect 3418 16028 3424 16040
rect 2823 16000 3424 16028
rect 2823 15997 2835 16000
rect 2777 15991 2835 15997
rect 3418 15988 3424 16000
rect 3476 15988 3482 16040
rect 3602 15988 3608 16040
rect 3660 16028 3666 16040
rect 3789 16031 3847 16037
rect 3789 16028 3801 16031
rect 3660 16000 3801 16028
rect 3660 15988 3666 16000
rect 3789 15997 3801 16000
rect 3835 15997 3847 16031
rect 3789 15991 3847 15997
rect 3878 15988 3884 16040
rect 3936 16028 3942 16040
rect 4065 16031 4123 16037
rect 4065 16028 4077 16031
rect 3936 16000 4077 16028
rect 3936 15988 3942 16000
rect 4065 15997 4077 16000
rect 4111 15997 4123 16031
rect 4065 15991 4123 15997
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 4801 16031 4859 16037
rect 4801 16028 4813 16031
rect 4396 16000 4813 16028
rect 4396 15988 4402 16000
rect 4801 15997 4813 16000
rect 4847 15997 4859 16031
rect 4801 15991 4859 15997
rect 5169 16031 5227 16037
rect 5169 15997 5181 16031
rect 5215 15997 5227 16031
rect 5169 15991 5227 15997
rect 5184 15960 5212 15991
rect 7926 15960 7932 15972
rect 5184 15932 7932 15960
rect 7926 15920 7932 15932
rect 7984 15920 7990 15972
rect 1397 15895 1455 15901
rect 1397 15861 1409 15895
rect 1443 15892 1455 15895
rect 2130 15892 2136 15904
rect 1443 15864 2136 15892
rect 1443 15861 1455 15864
rect 1397 15855 1455 15861
rect 2130 15852 2136 15864
rect 2188 15852 2194 15904
rect 3050 15852 3056 15904
rect 3108 15892 3114 15904
rect 5258 15892 5264 15904
rect 3108 15864 5264 15892
rect 3108 15852 3114 15864
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 5629 15895 5687 15901
rect 5629 15861 5641 15895
rect 5675 15892 5687 15895
rect 6086 15892 6092 15904
rect 5675 15864 6092 15892
rect 5675 15861 5687 15864
rect 5629 15855 5687 15861
rect 6086 15852 6092 15864
rect 6144 15852 6150 15904
rect 1104 15802 16836 15824
rect 1104 15750 2924 15802
rect 2976 15750 2988 15802
rect 3040 15750 3052 15802
rect 3104 15750 3116 15802
rect 3168 15750 3180 15802
rect 3232 15750 6872 15802
rect 6924 15750 6936 15802
rect 6988 15750 7000 15802
rect 7052 15750 7064 15802
rect 7116 15750 7128 15802
rect 7180 15750 10820 15802
rect 10872 15750 10884 15802
rect 10936 15750 10948 15802
rect 11000 15750 11012 15802
rect 11064 15750 11076 15802
rect 11128 15750 14768 15802
rect 14820 15750 14832 15802
rect 14884 15750 14896 15802
rect 14948 15750 14960 15802
rect 15012 15750 15024 15802
rect 15076 15750 16836 15802
rect 1104 15728 16836 15750
rect 4798 15648 4804 15700
rect 4856 15688 4862 15700
rect 5077 15691 5135 15697
rect 5077 15688 5089 15691
rect 4856 15660 5089 15688
rect 4856 15648 4862 15660
rect 5077 15657 5089 15660
rect 5123 15657 5135 15691
rect 5077 15651 5135 15657
rect 5258 15648 5264 15700
rect 5316 15688 5322 15700
rect 9582 15688 9588 15700
rect 5316 15660 9588 15688
rect 5316 15648 5322 15660
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 3145 15623 3203 15629
rect 3145 15589 3157 15623
rect 3191 15620 3203 15623
rect 6454 15620 6460 15632
rect 3191 15592 6460 15620
rect 3191 15589 3203 15592
rect 3145 15583 3203 15589
rect 6454 15580 6460 15592
rect 6512 15580 6518 15632
rect 4154 15512 4160 15564
rect 4212 15552 4218 15564
rect 5353 15555 5411 15561
rect 5353 15552 5365 15555
rect 4212 15524 5365 15552
rect 4212 15512 4218 15524
rect 5353 15521 5365 15524
rect 5399 15521 5411 15555
rect 5353 15515 5411 15521
rect 5445 15555 5503 15561
rect 5445 15521 5457 15555
rect 5491 15552 5503 15555
rect 5718 15552 5724 15564
rect 5491 15524 5724 15552
rect 5491 15521 5503 15524
rect 5445 15515 5503 15521
rect 5718 15512 5724 15524
rect 5776 15512 5782 15564
rect 1762 15484 1768 15496
rect 1723 15456 1768 15484
rect 1762 15444 1768 15456
rect 1820 15444 1826 15496
rect 4338 15484 4344 15496
rect 4299 15456 4344 15484
rect 4338 15444 4344 15456
rect 4396 15444 4402 15496
rect 4614 15484 4620 15496
rect 4575 15456 4620 15484
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15453 5319 15487
rect 5261 15447 5319 15453
rect 5537 15487 5595 15493
rect 5537 15453 5549 15487
rect 5583 15484 5595 15487
rect 6178 15484 6184 15496
rect 5583 15456 6184 15484
rect 5583 15453 5595 15456
rect 5537 15447 5595 15453
rect 2032 15419 2090 15425
rect 2032 15385 2044 15419
rect 2078 15416 2090 15419
rect 4062 15416 4068 15428
rect 2078 15388 4068 15416
rect 2078 15385 2090 15388
rect 2032 15379 2090 15385
rect 4062 15376 4068 15388
rect 4120 15376 4126 15428
rect 5277 15416 5305 15447
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15484 6331 15487
rect 7374 15484 7380 15496
rect 6319 15456 7380 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 7190 15416 7196 15428
rect 5277 15388 7196 15416
rect 3602 15308 3608 15360
rect 3660 15348 3666 15360
rect 5277 15348 5305 15388
rect 7190 15376 7196 15388
rect 7248 15376 7254 15428
rect 3660 15320 5305 15348
rect 3660 15308 3666 15320
rect 5810 15308 5816 15360
rect 5868 15348 5874 15360
rect 6089 15351 6147 15357
rect 6089 15348 6101 15351
rect 5868 15320 6101 15348
rect 5868 15308 5874 15320
rect 6089 15317 6101 15320
rect 6135 15317 6147 15351
rect 6089 15311 6147 15317
rect 1104 15258 16836 15280
rect 1104 15206 4898 15258
rect 4950 15206 4962 15258
rect 5014 15206 5026 15258
rect 5078 15206 5090 15258
rect 5142 15206 5154 15258
rect 5206 15206 8846 15258
rect 8898 15206 8910 15258
rect 8962 15206 8974 15258
rect 9026 15206 9038 15258
rect 9090 15206 9102 15258
rect 9154 15206 12794 15258
rect 12846 15206 12858 15258
rect 12910 15206 12922 15258
rect 12974 15206 12986 15258
rect 13038 15206 13050 15258
rect 13102 15206 16836 15258
rect 1104 15184 16836 15206
rect 5629 15147 5687 15153
rect 5629 15113 5641 15147
rect 5675 15144 5687 15147
rect 8478 15144 8484 15156
rect 5675 15116 8484 15144
rect 5675 15113 5687 15116
rect 5629 15107 5687 15113
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 3872 15079 3930 15085
rect 3872 15045 3884 15079
rect 3918 15076 3930 15079
rect 4062 15076 4068 15088
rect 3918 15048 4068 15076
rect 3918 15045 3930 15048
rect 3872 15039 3930 15045
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 6549 15079 6607 15085
rect 6549 15045 6561 15079
rect 6595 15076 6607 15079
rect 8570 15076 8576 15088
rect 6595 15048 8576 15076
rect 6595 15045 6607 15048
rect 6549 15039 6607 15045
rect 8570 15036 8576 15048
rect 8628 15036 8634 15088
rect 2032 15011 2090 15017
rect 2032 14977 2044 15011
rect 2078 15008 2090 15011
rect 4246 15008 4252 15020
rect 2078 14980 4252 15008
rect 2078 14977 2090 14980
rect 2032 14971 2090 14977
rect 4246 14968 4252 14980
rect 4304 14968 4310 15020
rect 5718 15008 5724 15020
rect 5679 14980 5724 15008
rect 5718 14968 5724 14980
rect 5776 14968 5782 15020
rect 5813 15011 5871 15017
rect 5813 14977 5825 15011
rect 5859 15008 5871 15011
rect 5994 15008 6000 15020
rect 5859 14980 6000 15008
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 5994 14968 6000 14980
rect 6052 14968 6058 15020
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 15008 6699 15011
rect 7006 15008 7012 15020
rect 6687 14980 7012 15008
rect 6687 14977 6699 14980
rect 6641 14971 6699 14977
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 3418 14900 3424 14952
rect 3476 14940 3482 14952
rect 3605 14943 3663 14949
rect 3605 14940 3617 14943
rect 3476 14912 3617 14940
rect 3476 14900 3482 14912
rect 3605 14909 3617 14912
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 5350 14900 5356 14952
rect 5408 14940 5414 14952
rect 5445 14943 5503 14949
rect 5445 14940 5457 14943
rect 5408 14912 5457 14940
rect 5408 14900 5414 14912
rect 5445 14909 5457 14912
rect 5491 14909 5503 14943
rect 6380 14940 6408 14971
rect 7006 14968 7012 14980
rect 7064 14968 7070 15020
rect 7098 14968 7104 15020
rect 7156 15008 7162 15020
rect 7156 14980 7201 15008
rect 7156 14968 7162 14980
rect 8754 14940 8760 14952
rect 6380 14912 8760 14940
rect 5445 14903 5503 14909
rect 8754 14900 8760 14912
rect 8812 14900 8818 14952
rect 6362 14872 6368 14884
rect 6323 14844 6368 14872
rect 6362 14832 6368 14844
rect 6420 14832 6426 14884
rect 7006 14832 7012 14884
rect 7064 14872 7070 14884
rect 8386 14872 8392 14884
rect 7064 14844 8392 14872
rect 7064 14832 7070 14844
rect 8386 14832 8392 14844
rect 8444 14832 8450 14884
rect 3145 14807 3203 14813
rect 3145 14773 3157 14807
rect 3191 14804 3203 14807
rect 4522 14804 4528 14816
rect 3191 14776 4528 14804
rect 3191 14773 3203 14776
rect 3145 14767 3203 14773
rect 4522 14764 4528 14776
rect 4580 14764 4586 14816
rect 4614 14764 4620 14816
rect 4672 14804 4678 14816
rect 4985 14807 5043 14813
rect 4985 14804 4997 14807
rect 4672 14776 4997 14804
rect 4672 14764 4678 14776
rect 4985 14773 4997 14776
rect 5031 14773 5043 14807
rect 5534 14804 5540 14816
rect 5495 14776 5540 14804
rect 4985 14767 5043 14773
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14804 7343 14807
rect 8294 14804 8300 14816
rect 7331 14776 8300 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 1104 14714 16836 14736
rect 1104 14662 2924 14714
rect 2976 14662 2988 14714
rect 3040 14662 3052 14714
rect 3104 14662 3116 14714
rect 3168 14662 3180 14714
rect 3232 14662 6872 14714
rect 6924 14662 6936 14714
rect 6988 14662 7000 14714
rect 7052 14662 7064 14714
rect 7116 14662 7128 14714
rect 7180 14662 10820 14714
rect 10872 14662 10884 14714
rect 10936 14662 10948 14714
rect 11000 14662 11012 14714
rect 11064 14662 11076 14714
rect 11128 14662 14768 14714
rect 14820 14662 14832 14714
rect 14884 14662 14896 14714
rect 14948 14662 14960 14714
rect 15012 14662 15024 14714
rect 15076 14662 16836 14714
rect 1104 14640 16836 14662
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14600 2835 14603
rect 4154 14600 4160 14612
rect 2823 14572 4160 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 4580 14572 6132 14600
rect 4580 14560 4586 14572
rect 5442 14492 5448 14544
rect 5500 14532 5506 14544
rect 5629 14535 5687 14541
rect 5629 14532 5641 14535
rect 5500 14504 5641 14532
rect 5500 14492 5506 14504
rect 5629 14501 5641 14504
rect 5675 14501 5687 14535
rect 5629 14495 5687 14501
rect 6104 14473 6132 14572
rect 6178 14560 6184 14612
rect 6236 14600 6242 14612
rect 6825 14603 6883 14609
rect 6825 14600 6837 14603
rect 6236 14572 6837 14600
rect 6236 14560 6242 14572
rect 6825 14569 6837 14572
rect 6871 14569 6883 14603
rect 6825 14563 6883 14569
rect 6546 14492 6552 14544
rect 6604 14532 6610 14544
rect 7929 14535 7987 14541
rect 7929 14532 7941 14535
rect 6604 14504 7941 14532
rect 6604 14492 6610 14504
rect 7929 14501 7941 14504
rect 7975 14501 7987 14535
rect 7929 14495 7987 14501
rect 6089 14467 6147 14473
rect 6089 14433 6101 14467
rect 6135 14433 6147 14467
rect 6089 14427 6147 14433
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14464 6331 14467
rect 6914 14464 6920 14476
rect 6319 14436 6920 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7190 14464 7196 14476
rect 7024 14436 7196 14464
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 2222 14396 2228 14408
rect 1443 14368 2228 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 1780 14340 1808 14368
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 7024 14405 7052 14436
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 9306 14464 9312 14476
rect 7484 14436 9312 14464
rect 5169 14399 5227 14405
rect 5169 14365 5181 14399
rect 5215 14396 5227 14399
rect 7009 14399 7067 14405
rect 5215 14368 6960 14396
rect 5215 14365 5227 14368
rect 5169 14359 5227 14365
rect 1670 14337 1676 14340
rect 1664 14328 1676 14337
rect 1631 14300 1676 14328
rect 1664 14291 1676 14300
rect 1670 14288 1676 14291
rect 1728 14288 1734 14340
rect 1762 14288 1768 14340
rect 1820 14288 1826 14340
rect 2038 14288 2044 14340
rect 2096 14328 2102 14340
rect 4430 14328 4436 14340
rect 2096 14300 4436 14328
rect 2096 14288 2102 14300
rect 4430 14288 4436 14300
rect 4488 14328 4494 14340
rect 4902 14331 4960 14337
rect 4902 14328 4914 14331
rect 4488 14300 4914 14328
rect 4488 14288 4494 14300
rect 4902 14297 4914 14300
rect 4948 14297 4960 14331
rect 6932 14328 6960 14368
rect 7009 14365 7021 14399
rect 7055 14365 7067 14399
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7009 14359 7067 14365
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7484 14405 7512 14436
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 7392 14368 7481 14396
rect 7190 14328 7196 14340
rect 6932 14300 7196 14328
rect 4902 14291 4960 14297
rect 3786 14260 3792 14272
rect 3747 14232 3792 14260
rect 3786 14220 3792 14232
rect 3844 14220 3850 14272
rect 4908 14260 4936 14291
rect 7190 14288 7196 14300
rect 7248 14288 7254 14340
rect 5810 14260 5816 14272
rect 4908 14232 5816 14260
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 5994 14260 6000 14272
rect 5955 14232 6000 14260
rect 5994 14220 6000 14232
rect 6052 14220 6058 14272
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 7392 14260 7420 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 8128 14328 8156 14359
rect 7484 14300 8156 14328
rect 7484 14272 7512 14300
rect 6420 14232 7420 14260
rect 6420 14220 6426 14232
rect 7466 14220 7472 14272
rect 7524 14220 7530 14272
rect 1104 14170 16836 14192
rect 1104 14118 4898 14170
rect 4950 14118 4962 14170
rect 5014 14118 5026 14170
rect 5078 14118 5090 14170
rect 5142 14118 5154 14170
rect 5206 14118 8846 14170
rect 8898 14118 8910 14170
rect 8962 14118 8974 14170
rect 9026 14118 9038 14170
rect 9090 14118 9102 14170
rect 9154 14118 12794 14170
rect 12846 14118 12858 14170
rect 12910 14118 12922 14170
rect 12974 14118 12986 14170
rect 13038 14118 13050 14170
rect 13102 14118 16836 14170
rect 1104 14096 16836 14118
rect 3145 14059 3203 14065
rect 3145 14025 3157 14059
rect 3191 14056 3203 14059
rect 6733 14059 6791 14065
rect 6733 14056 6745 14059
rect 3191 14028 6745 14056
rect 3191 14025 3203 14028
rect 3145 14019 3203 14025
rect 6733 14025 6745 14028
rect 6779 14025 6791 14059
rect 6733 14019 6791 14025
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 8481 14059 8539 14065
rect 8481 14056 8493 14059
rect 6880 14028 8493 14056
rect 6880 14016 6886 14028
rect 8481 14025 8493 14028
rect 8527 14025 8539 14059
rect 8481 14019 8539 14025
rect 3970 13988 3976 14000
rect 1780 13960 3976 13988
rect 1780 13929 1808 13960
rect 2038 13929 2044 13932
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13889 1823 13923
rect 2032 13920 2044 13929
rect 1999 13892 2044 13920
rect 1765 13883 1823 13889
rect 2032 13883 2044 13892
rect 2038 13880 2044 13883
rect 2096 13880 2102 13932
rect 3620 13929 3648 13960
rect 3970 13948 3976 13960
rect 4028 13948 4034 14000
rect 4062 13948 4068 14000
rect 4120 13948 4126 14000
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 3872 13923 3930 13929
rect 3872 13889 3884 13923
rect 3918 13920 3930 13923
rect 4080 13920 4108 13948
rect 5534 13920 5540 13932
rect 3918 13892 4108 13920
rect 5495 13892 5540 13920
rect 3918 13889 3930 13892
rect 3872 13883 3930 13889
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 5629 13923 5687 13929
rect 5629 13889 5641 13923
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5442 13852 5448 13864
rect 5000 13824 5448 13852
rect 5000 13793 5028 13824
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 4985 13787 5043 13793
rect 4985 13753 4997 13787
rect 5031 13753 5043 13787
rect 4985 13747 5043 13753
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 5442 13716 5448 13728
rect 1728 13688 5448 13716
rect 1728 13676 1734 13688
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 5644 13716 5672 13883
rect 5902 13880 5908 13932
rect 5960 13920 5966 13932
rect 7617 13923 7675 13929
rect 7617 13920 7629 13923
rect 5960 13892 7629 13920
rect 5960 13880 5966 13892
rect 7617 13889 7629 13892
rect 7663 13889 7675 13923
rect 7742 13920 7748 13932
rect 7703 13892 7748 13920
rect 7617 13883 7675 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 8202 13920 8208 13932
rect 7883 13892 8208 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 8662 13880 8668 13932
rect 8720 13920 8726 13932
rect 9309 13923 9367 13929
rect 8720 13892 8765 13920
rect 8720 13880 8726 13892
rect 9309 13889 9321 13923
rect 9355 13920 9367 13923
rect 11606 13920 11612 13932
rect 9355 13892 11612 13920
rect 9355 13889 9367 13892
rect 9309 13883 9367 13889
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 5718 13812 5724 13864
rect 5776 13852 5782 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 5776 13824 6837 13852
rect 5776 13812 5782 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 8018 13852 8024 13864
rect 6972 13824 7065 13852
rect 7116 13824 7696 13852
rect 7979 13824 8024 13852
rect 6972 13812 6978 13824
rect 5813 13787 5871 13793
rect 5813 13753 5825 13787
rect 5859 13784 5871 13787
rect 5902 13784 5908 13796
rect 5859 13756 5908 13784
rect 5859 13753 5871 13756
rect 5813 13747 5871 13753
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 6270 13744 6276 13796
rect 6328 13784 6334 13796
rect 6365 13787 6423 13793
rect 6365 13784 6377 13787
rect 6328 13756 6377 13784
rect 6328 13744 6334 13756
rect 6365 13753 6377 13756
rect 6411 13753 6423 13787
rect 6365 13747 6423 13753
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 6932 13784 6960 13812
rect 6788 13756 6960 13784
rect 6788 13744 6794 13756
rect 7116 13716 7144 13824
rect 7668 13784 7696 13824
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 9950 13852 9956 13864
rect 8404 13824 9956 13852
rect 8404 13784 8432 13824
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 7668 13756 8432 13784
rect 5644 13688 7144 13716
rect 7190 13676 7196 13728
rect 7248 13716 7254 13728
rect 9125 13719 9183 13725
rect 9125 13716 9137 13719
rect 7248 13688 9137 13716
rect 7248 13676 7254 13688
rect 9125 13685 9137 13688
rect 9171 13685 9183 13719
rect 9125 13679 9183 13685
rect 1104 13626 16836 13648
rect 1104 13574 2924 13626
rect 2976 13574 2988 13626
rect 3040 13574 3052 13626
rect 3104 13574 3116 13626
rect 3168 13574 3180 13626
rect 3232 13574 6872 13626
rect 6924 13574 6936 13626
rect 6988 13574 7000 13626
rect 7052 13574 7064 13626
rect 7116 13574 7128 13626
rect 7180 13574 10820 13626
rect 10872 13574 10884 13626
rect 10936 13574 10948 13626
rect 11000 13574 11012 13626
rect 11064 13574 11076 13626
rect 11128 13574 14768 13626
rect 14820 13574 14832 13626
rect 14884 13574 14896 13626
rect 14948 13574 14960 13626
rect 15012 13574 15024 13626
rect 15076 13574 16836 13626
rect 1104 13552 16836 13574
rect 3053 13515 3111 13521
rect 3053 13481 3065 13515
rect 3099 13512 3111 13515
rect 5169 13515 5227 13521
rect 3099 13484 5120 13512
rect 3099 13481 3111 13484
rect 3053 13475 3111 13481
rect 5092 13444 5120 13484
rect 5169 13481 5181 13515
rect 5215 13512 5227 13515
rect 5994 13512 6000 13524
rect 5215 13484 6000 13512
rect 5215 13481 5227 13484
rect 5169 13475 5227 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 7282 13512 7288 13524
rect 6104 13484 7288 13512
rect 6104 13444 6132 13484
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 9582 13472 9588 13524
rect 9640 13512 9646 13524
rect 11054 13512 11060 13524
rect 9640 13484 11060 13512
rect 9640 13472 9646 13484
rect 11054 13472 11060 13484
rect 11112 13472 11118 13524
rect 5092 13416 6132 13444
rect 7742 13404 7748 13456
rect 7800 13444 7806 13456
rect 9677 13447 9735 13453
rect 9677 13444 9689 13447
rect 7800 13416 9689 13444
rect 7800 13404 7806 13416
rect 9677 13413 9689 13416
rect 9723 13413 9735 13447
rect 9677 13407 9735 13413
rect 5442 13336 5448 13388
rect 5500 13376 5506 13388
rect 7929 13379 7987 13385
rect 7929 13376 7941 13379
rect 5500 13348 5948 13376
rect 5500 13336 5506 13348
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 1719 13280 3801 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 3789 13277 3801 13280
rect 3835 13308 3847 13311
rect 3878 13308 3884 13320
rect 3835 13280 3884 13308
rect 3835 13277 3847 13280
rect 3789 13271 3847 13277
rect 3878 13268 3884 13280
rect 3936 13268 3942 13320
rect 3988 13280 5764 13308
rect 1762 13200 1768 13252
rect 1820 13240 1826 13252
rect 1918 13243 1976 13249
rect 1918 13240 1930 13243
rect 1820 13212 1930 13240
rect 1820 13200 1826 13212
rect 1918 13209 1930 13212
rect 1964 13209 1976 13243
rect 1918 13203 1976 13209
rect 2038 13200 2044 13252
rect 2096 13240 2102 13252
rect 3988 13240 4016 13280
rect 2096 13212 4016 13240
rect 4056 13243 4114 13249
rect 2096 13200 2102 13212
rect 4056 13209 4068 13243
rect 4102 13240 4114 13243
rect 4246 13240 4252 13252
rect 4102 13212 4252 13240
rect 4102 13209 4114 13212
rect 4056 13203 4114 13209
rect 4246 13200 4252 13212
rect 4304 13200 4310 13252
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 5629 13175 5687 13181
rect 5629 13172 5641 13175
rect 3384 13144 5641 13172
rect 3384 13132 3390 13144
rect 5629 13141 5641 13144
rect 5675 13141 5687 13175
rect 5736 13172 5764 13280
rect 5920 13240 5948 13348
rect 6932 13348 7941 13376
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 6932 13308 6960 13348
rect 7929 13345 7941 13348
rect 7975 13345 7987 13379
rect 7929 13339 7987 13345
rect 8021 13379 8079 13385
rect 8021 13345 8033 13379
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 6512 13280 6960 13308
rect 7009 13311 7067 13317
rect 6512 13268 6518 13280
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 7190 13308 7196 13320
rect 7055 13280 7196 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 7558 13268 7564 13320
rect 7616 13308 7622 13320
rect 7837 13311 7895 13317
rect 7837 13308 7849 13311
rect 7616 13280 7849 13308
rect 7616 13268 7622 13280
rect 7837 13277 7849 13280
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 6086 13240 6092 13252
rect 5920 13212 6092 13240
rect 6086 13200 6092 13212
rect 6144 13240 6150 13252
rect 6546 13240 6552 13252
rect 6144 13212 6552 13240
rect 6144 13200 6150 13212
rect 6546 13200 6552 13212
rect 6604 13240 6610 13252
rect 6742 13243 6800 13249
rect 6742 13240 6754 13243
rect 6604 13212 6754 13240
rect 6604 13200 6610 13212
rect 6742 13209 6754 13212
rect 6788 13209 6800 13243
rect 6742 13203 6800 13209
rect 6914 13200 6920 13252
rect 6972 13240 6978 13252
rect 7282 13240 7288 13252
rect 6972 13212 7288 13240
rect 6972 13200 6978 13212
rect 7282 13200 7288 13212
rect 7340 13240 7346 13252
rect 8036 13240 8064 13339
rect 8754 13336 8760 13388
rect 8812 13376 8818 13388
rect 9033 13379 9091 13385
rect 9033 13376 9045 13379
rect 8812 13348 9045 13376
rect 8812 13336 8818 13348
rect 9033 13345 9045 13348
rect 9079 13376 9091 13379
rect 10686 13376 10692 13388
rect 9079 13348 10692 13376
rect 9079 13345 9091 13348
rect 9033 13339 9091 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 8386 13268 8392 13320
rect 8444 13308 8450 13320
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 8444 13280 8953 13308
rect 8444 13268 8450 13280
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 9858 13308 9864 13320
rect 9819 13280 9864 13308
rect 8941 13271 8999 13277
rect 7340 13212 8064 13240
rect 8956 13240 8984 13271
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 9217 13243 9275 13249
rect 8956 13212 9076 13240
rect 7340 13200 7346 13212
rect 7469 13175 7527 13181
rect 7469 13172 7481 13175
rect 5736 13144 7481 13172
rect 5629 13135 5687 13141
rect 7469 13141 7481 13144
rect 7515 13141 7527 13175
rect 7469 13135 7527 13141
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8941 13175 8999 13181
rect 8941 13172 8953 13175
rect 8076 13144 8953 13172
rect 8076 13132 8082 13144
rect 8941 13141 8953 13144
rect 8987 13141 8999 13175
rect 9048 13172 9076 13212
rect 9217 13209 9229 13243
rect 9263 13240 9275 13243
rect 10502 13240 10508 13252
rect 9263 13212 10508 13240
rect 9263 13209 9275 13212
rect 9217 13203 9275 13209
rect 10502 13200 10508 13212
rect 10560 13200 10566 13252
rect 11238 13172 11244 13184
rect 9048 13144 11244 13172
rect 8941 13135 8999 13141
rect 11238 13132 11244 13144
rect 11296 13132 11302 13184
rect 1104 13082 16836 13104
rect 1104 13030 4898 13082
rect 4950 13030 4962 13082
rect 5014 13030 5026 13082
rect 5078 13030 5090 13082
rect 5142 13030 5154 13082
rect 5206 13030 8846 13082
rect 8898 13030 8910 13082
rect 8962 13030 8974 13082
rect 9026 13030 9038 13082
rect 9090 13030 9102 13082
rect 9154 13030 12794 13082
rect 12846 13030 12858 13082
rect 12910 13030 12922 13082
rect 12974 13030 12986 13082
rect 13038 13030 13050 13082
rect 13102 13030 16836 13082
rect 1104 13008 16836 13030
rect 1394 12968 1400 12980
rect 1355 12940 1400 12968
rect 1394 12928 1400 12940
rect 1452 12928 1458 12980
rect 2222 12928 2228 12980
rect 2280 12968 2286 12980
rect 5718 12968 5724 12980
rect 2280 12940 4384 12968
rect 5679 12940 5724 12968
rect 2280 12928 2286 12940
rect 4356 12900 4384 12940
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 6546 12928 6552 12980
rect 6604 12968 6610 12980
rect 8294 12968 8300 12980
rect 6604 12940 8300 12968
rect 6604 12928 6610 12940
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 11974 12968 11980 12980
rect 9324 12940 11980 12968
rect 8018 12900 8024 12912
rect 4356 12872 8024 12900
rect 1578 12832 1584 12844
rect 1539 12804 1584 12832
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 2682 12792 2688 12844
rect 2740 12832 2746 12844
rect 2958 12832 2964 12844
rect 2740 12804 2785 12832
rect 2919 12804 2964 12832
rect 2740 12792 2746 12804
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3786 12792 3792 12844
rect 3844 12832 3850 12844
rect 4356 12841 4384 12872
rect 8018 12860 8024 12872
rect 8076 12860 8082 12912
rect 8665 12903 8723 12909
rect 8665 12869 8677 12903
rect 8711 12900 8723 12903
rect 9030 12900 9036 12912
rect 8711 12872 9036 12900
rect 8711 12869 8723 12872
rect 8665 12863 8723 12869
rect 9030 12860 9036 12872
rect 9088 12860 9094 12912
rect 9324 12909 9352 12940
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 9309 12903 9367 12909
rect 9309 12869 9321 12903
rect 9355 12869 9367 12903
rect 9309 12863 9367 12869
rect 3881 12835 3939 12841
rect 3881 12832 3893 12835
rect 3844 12804 3893 12832
rect 3844 12792 3850 12804
rect 3881 12801 3893 12804
rect 3927 12801 3939 12835
rect 3881 12795 3939 12801
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 4430 12792 4436 12844
rect 4488 12832 4494 12844
rect 4608 12835 4666 12841
rect 4608 12832 4620 12835
rect 4488 12804 4620 12832
rect 4488 12792 4494 12804
rect 4608 12801 4620 12804
rect 4654 12832 4666 12835
rect 7478 12835 7536 12841
rect 7478 12832 7490 12835
rect 4654 12804 7490 12832
rect 4654 12801 4666 12804
rect 4608 12795 4666 12801
rect 7478 12801 7490 12804
rect 7524 12801 7536 12835
rect 7478 12795 7536 12801
rect 7650 12792 7656 12844
rect 7708 12832 7714 12844
rect 7745 12835 7803 12841
rect 7745 12832 7757 12835
rect 7708 12804 7757 12832
rect 7708 12792 7714 12804
rect 7745 12801 7757 12804
rect 7791 12832 7803 12835
rect 8389 12835 8447 12841
rect 7791 12804 8064 12832
rect 7791 12801 7803 12804
rect 7745 12795 7803 12801
rect 8036 12776 8064 12804
rect 8389 12801 8401 12835
rect 8435 12832 8447 12835
rect 8846 12832 8852 12844
rect 8435 12804 8852 12832
rect 8435 12801 8447 12804
rect 8389 12795 8447 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9953 12835 10011 12841
rect 9539 12804 9904 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 2041 12767 2099 12773
rect 2041 12733 2053 12767
rect 2087 12764 2099 12767
rect 2314 12764 2320 12776
rect 2087 12736 2320 12764
rect 2087 12733 2099 12736
rect 2041 12727 2099 12733
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 2844 12767 2902 12773
rect 2844 12733 2856 12767
rect 2890 12764 2902 12767
rect 3697 12767 3755 12773
rect 2890 12736 3648 12764
rect 2890 12733 2902 12736
rect 2844 12727 2902 12733
rect 3237 12699 3295 12705
rect 3237 12665 3249 12699
rect 3283 12696 3295 12699
rect 3418 12696 3424 12708
rect 3283 12668 3424 12696
rect 3283 12665 3295 12668
rect 3237 12659 3295 12665
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 3620 12628 3648 12736
rect 3697 12733 3709 12767
rect 3743 12764 3755 12767
rect 4154 12764 4160 12776
rect 3743 12736 4160 12764
rect 3743 12733 3755 12736
rect 3697 12727 3755 12733
rect 4154 12724 4160 12736
rect 4212 12724 4218 12776
rect 8018 12724 8024 12776
rect 8076 12724 8082 12776
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12764 8631 12767
rect 9674 12764 9680 12776
rect 8619 12736 9680 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 8938 12656 8944 12708
rect 8996 12696 9002 12708
rect 9125 12699 9183 12705
rect 9125 12696 9137 12699
rect 8996 12668 9137 12696
rect 8996 12656 9002 12668
rect 9125 12665 9137 12668
rect 9171 12665 9183 12699
rect 9125 12659 9183 12665
rect 9876 12696 9904 12804
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10042 12832 10048 12844
rect 9999 12804 10048 12832
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12832 10655 12835
rect 11054 12832 11060 12844
rect 10643 12804 11060 12832
rect 10643 12801 10655 12804
rect 10597 12795 10655 12801
rect 11054 12792 11060 12804
rect 11112 12832 11118 12844
rect 11422 12832 11428 12844
rect 11112 12804 11428 12832
rect 11112 12792 11118 12804
rect 11422 12792 11428 12804
rect 11480 12792 11486 12844
rect 12158 12696 12164 12708
rect 9876 12668 12164 12696
rect 6365 12631 6423 12637
rect 6365 12628 6377 12631
rect 3620 12600 6377 12628
rect 6365 12597 6377 12600
rect 6411 12597 6423 12631
rect 6365 12591 6423 12597
rect 7742 12588 7748 12640
rect 7800 12628 7806 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 7800 12600 8217 12628
rect 7800 12588 7806 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8386 12628 8392 12640
rect 8347 12600 8392 12628
rect 8205 12591 8263 12597
rect 8386 12588 8392 12600
rect 8444 12588 8450 12640
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 9214 12628 9220 12640
rect 8536 12600 9220 12628
rect 8536 12588 8542 12600
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 9490 12588 9496 12640
rect 9548 12628 9554 12640
rect 9876 12628 9904 12668
rect 12158 12656 12164 12668
rect 12216 12656 12222 12708
rect 9548 12600 9904 12628
rect 10045 12631 10103 12637
rect 9548 12588 9554 12600
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10134 12628 10140 12640
rect 10091 12600 10140 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 10226 12588 10232 12640
rect 10284 12628 10290 12640
rect 10781 12631 10839 12637
rect 10781 12628 10793 12631
rect 10284 12600 10793 12628
rect 10284 12588 10290 12600
rect 10781 12597 10793 12600
rect 10827 12597 10839 12631
rect 10781 12591 10839 12597
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 12066 12628 12072 12640
rect 11296 12600 12072 12628
rect 11296 12588 11302 12600
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 1104 12538 16836 12560
rect 1104 12486 2924 12538
rect 2976 12486 2988 12538
rect 3040 12486 3052 12538
rect 3104 12486 3116 12538
rect 3168 12486 3180 12538
rect 3232 12486 6872 12538
rect 6924 12486 6936 12538
rect 6988 12486 7000 12538
rect 7052 12486 7064 12538
rect 7116 12486 7128 12538
rect 7180 12486 10820 12538
rect 10872 12486 10884 12538
rect 10936 12486 10948 12538
rect 11000 12486 11012 12538
rect 11064 12486 11076 12538
rect 11128 12486 14768 12538
rect 14820 12486 14832 12538
rect 14884 12486 14896 12538
rect 14948 12486 14960 12538
rect 15012 12486 15024 12538
rect 15076 12486 16836 12538
rect 1104 12464 16836 12486
rect 1397 12427 1455 12433
rect 1397 12393 1409 12427
rect 1443 12424 1455 12427
rect 2774 12424 2780 12436
rect 1443 12396 2780 12424
rect 1443 12393 1455 12396
rect 1397 12387 1455 12393
rect 2774 12384 2780 12396
rect 2832 12384 2838 12436
rect 3970 12384 3976 12436
rect 4028 12424 4034 12436
rect 7650 12424 7656 12436
rect 4028 12396 7656 12424
rect 4028 12384 4034 12396
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 7926 12424 7932 12436
rect 7887 12396 7932 12424
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 8294 12424 8300 12436
rect 8255 12396 8300 12424
rect 8294 12384 8300 12396
rect 8352 12424 8358 12436
rect 10410 12424 10416 12436
rect 8352 12396 10416 12424
rect 8352 12384 8358 12396
rect 10410 12384 10416 12396
rect 10468 12424 10474 12436
rect 10778 12424 10784 12436
rect 10468 12396 10640 12424
rect 10739 12396 10784 12424
rect 10468 12384 10474 12396
rect 2593 12359 2651 12365
rect 2593 12325 2605 12359
rect 2639 12356 2651 12359
rect 3050 12356 3056 12368
rect 2639 12328 3056 12356
rect 2639 12325 2651 12328
rect 2593 12319 2651 12325
rect 3050 12316 3056 12328
rect 3108 12356 3114 12368
rect 3418 12356 3424 12368
rect 3108 12328 3424 12356
rect 3108 12316 3114 12328
rect 3418 12316 3424 12328
rect 3476 12316 3482 12368
rect 6089 12359 6147 12365
rect 6089 12356 6101 12359
rect 5460 12328 6101 12356
rect 2130 12248 2136 12300
rect 2188 12297 2194 12300
rect 2188 12291 2237 12297
rect 2188 12257 2191 12291
rect 2225 12257 2237 12291
rect 2188 12251 2237 12257
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 2498 12288 2504 12300
rect 2363 12260 2504 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2188 12248 2194 12251
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 3237 12291 3295 12297
rect 3237 12257 3249 12291
rect 3283 12288 3295 12291
rect 3326 12288 3332 12300
rect 3283 12260 3332 12288
rect 3283 12257 3295 12260
rect 3237 12251 3295 12257
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 4614 12297 4620 12300
rect 4433 12291 4491 12297
rect 4433 12288 4445 12291
rect 3896 12260 4445 12288
rect 2038 12180 2044 12232
rect 2096 12220 2102 12232
rect 3053 12223 3111 12229
rect 2096 12192 2141 12220
rect 2096 12180 2102 12192
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3786 12220 3792 12232
rect 3099 12192 3792 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3786 12180 3792 12192
rect 3844 12180 3850 12232
rect 3896 12152 3924 12260
rect 4433 12257 4445 12260
rect 4479 12257 4491 12291
rect 4433 12251 4491 12257
rect 4592 12291 4620 12297
rect 4592 12257 4604 12291
rect 4592 12251 4620 12257
rect 4614 12248 4620 12251
rect 4672 12248 4678 12300
rect 4982 12288 4988 12300
rect 4895 12260 4988 12288
rect 4982 12248 4988 12260
rect 5040 12288 5046 12300
rect 5460 12297 5488 12328
rect 6089 12325 6101 12328
rect 6135 12325 6147 12359
rect 6089 12319 6147 12325
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 8941 12359 8999 12365
rect 8941 12356 8953 12359
rect 8260 12328 8953 12356
rect 8260 12316 8266 12328
rect 8941 12325 8953 12328
rect 8987 12325 8999 12359
rect 10612 12356 10640 12396
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 11330 12424 11336 12436
rect 11291 12396 11336 12424
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 12066 12424 12072 12436
rect 12027 12396 12072 12424
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 12342 12356 12348 12368
rect 8941 12319 8999 12325
rect 9968 12328 10180 12356
rect 10612 12328 12348 12356
rect 5445 12291 5503 12297
rect 5040 12260 5304 12288
rect 5040 12248 5046 12260
rect 4706 12220 4712 12232
rect 4667 12192 4712 12220
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 5276 12220 5304 12260
rect 5445 12257 5457 12291
rect 5491 12257 5503 12291
rect 9968 12288 9996 12328
rect 5445 12251 5503 12257
rect 8956 12260 9996 12288
rect 8956 12232 8984 12260
rect 5626 12220 5632 12232
rect 5276 12192 5488 12220
rect 5587 12192 5632 12220
rect 3712 12124 3924 12152
rect 5460 12152 5488 12192
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 6178 12180 6184 12232
rect 6236 12220 6242 12232
rect 7469 12223 7527 12229
rect 7469 12220 7481 12223
rect 6236 12192 7481 12220
rect 6236 12180 6242 12192
rect 7469 12189 7481 12192
rect 7515 12189 7527 12223
rect 8110 12220 8116 12232
rect 8071 12192 8116 12220
rect 7469 12183 7527 12189
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12189 8263 12223
rect 8938 12220 8944 12232
rect 8205 12183 8263 12189
rect 8588 12192 8944 12220
rect 6362 12152 6368 12164
rect 5460 12124 6368 12152
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 3602 12084 3608 12096
rect 2096 12056 3608 12084
rect 2096 12044 2102 12056
rect 3602 12044 3608 12056
rect 3660 12084 3666 12096
rect 3712 12084 3740 12124
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 6454 12112 6460 12164
rect 6512 12152 6518 12164
rect 7224 12155 7282 12161
rect 6512 12124 7144 12152
rect 6512 12112 6518 12124
rect 3660 12056 3740 12084
rect 3789 12087 3847 12093
rect 3660 12044 3666 12056
rect 3789 12053 3801 12087
rect 3835 12084 3847 12087
rect 6822 12084 6828 12096
rect 3835 12056 6828 12084
rect 3835 12053 3847 12056
rect 3789 12047 3847 12053
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 7116 12084 7144 12124
rect 7224 12121 7236 12155
rect 7270 12152 7282 12155
rect 7650 12152 7656 12164
rect 7270 12124 7656 12152
rect 7270 12121 7282 12124
rect 7224 12115 7282 12121
rect 7650 12112 7656 12124
rect 7708 12112 7714 12164
rect 8220 12152 8248 12183
rect 8588 12164 8616 12192
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9122 12220 9128 12232
rect 9083 12192 9128 12220
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 9398 12220 9404 12232
rect 9355 12192 9404 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 8128 12124 8248 12152
rect 8389 12155 8447 12161
rect 8128 12096 8156 12124
rect 8389 12121 8401 12155
rect 8435 12152 8447 12155
rect 8570 12152 8576 12164
rect 8435 12124 8576 12152
rect 8435 12121 8447 12124
rect 8389 12115 8447 12121
rect 8570 12112 8576 12124
rect 8628 12112 8634 12164
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 9030 12152 9036 12164
rect 8720 12124 9036 12152
rect 8720 12112 8726 12124
rect 9030 12112 9036 12124
rect 9088 12112 9094 12164
rect 9240 12152 9268 12183
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 10042 12220 10048 12232
rect 10003 12192 10048 12220
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10152 12220 10180 12328
rect 12342 12316 12348 12328
rect 12400 12316 12406 12368
rect 10686 12288 10692 12300
rect 10647 12260 10692 12288
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 10597 12223 10655 12229
rect 10597 12220 10609 12223
rect 10152 12192 10609 12220
rect 10597 12189 10609 12192
rect 10643 12189 10655 12223
rect 11514 12220 11520 12232
rect 11475 12192 11520 12220
rect 10597 12183 10655 12189
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 11974 12220 11980 12232
rect 11935 12192 11980 12220
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 12158 12220 12164 12232
rect 12119 12192 12164 12220
rect 12158 12180 12164 12192
rect 12216 12180 12222 12232
rect 9240 12124 10088 12152
rect 8110 12084 8116 12096
rect 7116 12056 8116 12084
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 9953 12087 10011 12093
rect 9953 12084 9965 12087
rect 9732 12056 9965 12084
rect 9732 12044 9738 12056
rect 9953 12053 9965 12056
rect 9999 12053 10011 12087
rect 10060 12084 10088 12124
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 10778 12152 10784 12164
rect 10560 12124 10784 12152
rect 10560 12112 10566 12124
rect 10778 12112 10784 12124
rect 10836 12152 10842 12164
rect 10873 12155 10931 12161
rect 10873 12152 10885 12155
rect 10836 12124 10885 12152
rect 10836 12112 10842 12124
rect 10873 12121 10885 12124
rect 10919 12121 10931 12155
rect 10873 12115 10931 12121
rect 10134 12084 10140 12096
rect 10060 12056 10140 12084
rect 9953 12047 10011 12053
rect 10134 12044 10140 12056
rect 10192 12084 10198 12096
rect 11146 12084 11152 12096
rect 10192 12056 11152 12084
rect 10192 12044 10198 12056
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 1104 11994 16836 12016
rect 1104 11942 4898 11994
rect 4950 11942 4962 11994
rect 5014 11942 5026 11994
rect 5078 11942 5090 11994
rect 5142 11942 5154 11994
rect 5206 11942 8846 11994
rect 8898 11942 8910 11994
rect 8962 11942 8974 11994
rect 9026 11942 9038 11994
rect 9090 11942 9102 11994
rect 9154 11942 12794 11994
rect 12846 11942 12858 11994
rect 12910 11942 12922 11994
rect 12974 11942 12986 11994
rect 13038 11942 13050 11994
rect 13102 11942 16836 11994
rect 1104 11920 16836 11942
rect 1578 11840 1584 11892
rect 1636 11880 1642 11892
rect 1857 11883 1915 11889
rect 1857 11880 1869 11883
rect 1636 11852 1869 11880
rect 1636 11840 1642 11852
rect 1857 11849 1869 11852
rect 1903 11849 1915 11883
rect 4154 11880 4160 11892
rect 4115 11852 4160 11880
rect 1857 11843 1915 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5902 11840 5908 11892
rect 5960 11880 5966 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 5960 11852 8217 11880
rect 5960 11840 5966 11852
rect 8205 11849 8217 11852
rect 8251 11849 8263 11883
rect 8205 11843 8263 11849
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 10134 11880 10140 11892
rect 8628 11852 10140 11880
rect 8628 11840 8634 11852
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 4430 11772 4436 11824
rect 4488 11812 4494 11824
rect 5270 11815 5328 11821
rect 5270 11812 5282 11815
rect 4488 11784 5282 11812
rect 4488 11772 4494 11784
rect 5270 11781 5282 11784
rect 5316 11781 5328 11815
rect 5270 11775 5328 11781
rect 6638 11772 6644 11824
rect 6696 11812 6702 11824
rect 8294 11812 8300 11824
rect 6696 11784 8300 11812
rect 6696 11772 6702 11784
rect 8294 11772 8300 11784
rect 8352 11812 8358 11824
rect 10321 11815 10379 11821
rect 10321 11812 10333 11815
rect 8352 11784 8616 11812
rect 8352 11772 8358 11784
rect 5442 11704 5448 11756
rect 5500 11744 5506 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5500 11716 5549 11744
rect 5500 11704 5506 11716
rect 5537 11713 5549 11716
rect 5583 11744 5595 11747
rect 6178 11744 6184 11756
rect 5583 11716 6184 11744
rect 5583 11713 5595 11716
rect 5537 11707 5595 11713
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 7466 11704 7472 11756
rect 7524 11753 7530 11756
rect 7524 11744 7536 11753
rect 7745 11747 7803 11753
rect 7524 11716 7569 11744
rect 7524 11707 7536 11716
rect 7745 11713 7757 11747
rect 7791 11744 7803 11747
rect 8018 11744 8024 11756
rect 7791 11716 8024 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 7524 11704 7530 11707
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8588 11753 8616 11784
rect 9232 11784 10333 11812
rect 8573 11747 8631 11753
rect 8573 11713 8585 11747
rect 8619 11713 8631 11747
rect 8573 11707 8631 11713
rect 9030 11704 9036 11756
rect 9088 11744 9094 11756
rect 9232 11744 9260 11784
rect 10321 11781 10333 11784
rect 10367 11781 10379 11815
rect 10321 11775 10379 11781
rect 9088 11716 9260 11744
rect 9088 11704 9094 11716
rect 9398 11704 9404 11756
rect 9456 11744 9462 11756
rect 9493 11747 9551 11753
rect 9493 11744 9505 11747
rect 9456 11716 9505 11744
rect 9456 11704 9462 11716
rect 9493 11713 9505 11716
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 10192 11716 10517 11744
rect 10192 11704 10198 11716
rect 10505 11713 10517 11716
rect 10551 11744 10563 11747
rect 11330 11744 11336 11756
rect 10551 11716 11336 11744
rect 10551 11713 10563 11716
rect 10505 11707 10563 11713
rect 11330 11704 11336 11716
rect 11388 11704 11394 11756
rect 11698 11744 11704 11756
rect 11659 11716 11704 11744
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11713 12219 11747
rect 12342 11744 12348 11756
rect 12303 11716 12348 11744
rect 12161 11707 12219 11713
rect 2130 11636 2136 11688
rect 2188 11676 2194 11688
rect 2682 11685 2688 11688
rect 2501 11679 2559 11685
rect 2501 11676 2513 11679
rect 2188 11648 2513 11676
rect 2188 11636 2194 11648
rect 2501 11645 2513 11648
rect 2547 11645 2559 11679
rect 2501 11639 2559 11645
rect 2660 11679 2688 11685
rect 2660 11645 2672 11679
rect 2660 11639 2688 11645
rect 2682 11636 2688 11639
rect 2740 11636 2746 11688
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 3510 11676 3516 11688
rect 2832 11648 2877 11676
rect 3471 11648 3516 11676
rect 2832 11636 2838 11648
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 3694 11676 3700 11688
rect 3655 11648 3700 11676
rect 3694 11636 3700 11648
rect 3752 11636 3758 11688
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 8260 11648 8677 11676
rect 8260 11636 8266 11648
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 8938 11636 8944 11688
rect 8996 11676 9002 11688
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 8996 11648 9597 11676
rect 8996 11636 9002 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 3050 11608 3056 11620
rect 3011 11580 3056 11608
rect 3050 11568 3056 11580
rect 3108 11568 3114 11620
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 5810 11608 5816 11620
rect 5592 11580 5816 11608
rect 5592 11568 5598 11580
rect 5810 11568 5816 11580
rect 5868 11608 5874 11620
rect 9692 11608 9720 11639
rect 9766 11636 9772 11688
rect 9824 11676 9830 11688
rect 9824 11648 9869 11676
rect 9824 11636 9830 11648
rect 10226 11636 10232 11688
rect 10284 11676 10290 11688
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10284 11648 10793 11676
rect 10284 11636 10290 11648
rect 10781 11645 10793 11648
rect 10827 11676 10839 11679
rect 12176 11676 12204 11707
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 10827 11648 12204 11676
rect 10827 11645 10839 11648
rect 10781 11639 10839 11645
rect 11606 11608 11612 11620
rect 5868 11580 6500 11608
rect 5868 11568 5874 11580
rect 2682 11500 2688 11552
rect 2740 11540 2746 11552
rect 6365 11543 6423 11549
rect 6365 11540 6377 11543
rect 2740 11512 6377 11540
rect 2740 11500 2746 11512
rect 6365 11509 6377 11512
rect 6411 11509 6423 11543
rect 6472 11540 6500 11580
rect 8312 11580 9444 11608
rect 9692 11580 11612 11608
rect 7466 11540 7472 11552
rect 6472 11512 7472 11540
rect 6365 11503 6423 11509
rect 7466 11500 7472 11512
rect 7524 11540 7530 11552
rect 8312 11540 8340 11580
rect 7524 11512 8340 11540
rect 7524 11500 7530 11512
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 8849 11543 8907 11549
rect 8849 11540 8861 11543
rect 8812 11512 8861 11540
rect 8812 11500 8818 11512
rect 8849 11509 8861 11512
rect 8895 11540 8907 11543
rect 8938 11540 8944 11552
rect 8895 11512 8944 11540
rect 8895 11509 8907 11512
rect 8849 11503 8907 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9306 11540 9312 11552
rect 9267 11512 9312 11540
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9416 11540 9444 11580
rect 11606 11568 11612 11580
rect 11664 11568 11670 11620
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 9416 11512 10701 11540
rect 10689 11509 10701 11512
rect 10735 11540 10747 11543
rect 11517 11543 11575 11549
rect 11517 11540 11529 11543
rect 10735 11512 11529 11540
rect 10735 11509 10747 11512
rect 10689 11503 10747 11509
rect 11517 11509 11529 11512
rect 11563 11509 11575 11543
rect 11517 11503 11575 11509
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 12253 11543 12311 11549
rect 12253 11540 12265 11543
rect 11848 11512 12265 11540
rect 11848 11500 11854 11512
rect 12253 11509 12265 11512
rect 12299 11509 12311 11543
rect 12253 11503 12311 11509
rect 1104 11450 16836 11472
rect 1104 11398 2924 11450
rect 2976 11398 2988 11450
rect 3040 11398 3052 11450
rect 3104 11398 3116 11450
rect 3168 11398 3180 11450
rect 3232 11398 6872 11450
rect 6924 11398 6936 11450
rect 6988 11398 7000 11450
rect 7052 11398 7064 11450
rect 7116 11398 7128 11450
rect 7180 11398 10820 11450
rect 10872 11398 10884 11450
rect 10936 11398 10948 11450
rect 11000 11398 11012 11450
rect 11064 11398 11076 11450
rect 11128 11398 14768 11450
rect 14820 11398 14832 11450
rect 14884 11398 14896 11450
rect 14948 11398 14960 11450
rect 15012 11398 15024 11450
rect 15076 11398 16836 11450
rect 1104 11376 16836 11398
rect 1443 11339 1501 11345
rect 1443 11305 1455 11339
rect 1489 11336 1501 11339
rect 3786 11336 3792 11348
rect 1489 11308 3648 11336
rect 3747 11308 3792 11336
rect 1489 11305 1501 11308
rect 1443 11299 1501 11305
rect 3620 11268 3648 11308
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 4264 11308 5534 11336
rect 4264 11268 4292 11308
rect 3620 11240 4292 11268
rect 5506 11268 5534 11308
rect 5626 11296 5632 11348
rect 5684 11336 5690 11348
rect 5684 11308 5729 11336
rect 6104 11308 7328 11336
rect 5684 11296 5690 11308
rect 6104 11268 6132 11308
rect 5506 11240 6132 11268
rect 7300 11268 7328 11308
rect 7374 11296 7380 11348
rect 7432 11336 7438 11348
rect 7469 11339 7527 11345
rect 7469 11336 7481 11339
rect 7432 11308 7481 11336
rect 7432 11296 7438 11308
rect 7469 11305 7481 11308
rect 7515 11305 7527 11339
rect 7469 11299 7527 11305
rect 9677 11339 9735 11345
rect 9677 11305 9689 11339
rect 9723 11336 9735 11339
rect 9858 11336 9864 11348
rect 9723 11308 9864 11336
rect 9723 11305 9735 11308
rect 9677 11299 9735 11305
rect 9858 11296 9864 11308
rect 9916 11296 9922 11348
rect 9950 11296 9956 11348
rect 10008 11336 10014 11348
rect 10137 11339 10195 11345
rect 10137 11336 10149 11339
rect 10008 11308 10149 11336
rect 10008 11296 10014 11308
rect 10137 11305 10149 11308
rect 10183 11305 10195 11339
rect 10137 11299 10195 11305
rect 10318 11296 10324 11348
rect 10376 11336 10382 11348
rect 10778 11336 10784 11348
rect 10376 11308 10784 11336
rect 10376 11296 10382 11308
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 11606 11336 11612 11348
rect 11567 11308 11612 11336
rect 11606 11296 11612 11308
rect 11664 11336 11670 11348
rect 12618 11336 12624 11348
rect 11664 11308 12624 11336
rect 11664 11296 11670 11308
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 10042 11268 10048 11280
rect 7300 11240 10048 11268
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 10502 11228 10508 11280
rect 10560 11268 10566 11280
rect 13357 11271 13415 11277
rect 13357 11268 13369 11271
rect 10560 11240 13369 11268
rect 10560 11228 10566 11240
rect 13357 11237 13369 11240
rect 13403 11237 13415 11271
rect 13357 11231 13415 11237
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11200 2927 11203
rect 5169 11203 5227 11209
rect 2915 11172 4200 11200
rect 2915 11169 2927 11172
rect 2869 11163 2927 11169
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3418 11132 3424 11144
rect 3283 11104 3424 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 4172 11132 4200 11172
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 5442 11200 5448 11212
rect 5215 11172 5448 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 8018 11200 8024 11212
rect 7979 11172 8024 11200
rect 8018 11160 8024 11172
rect 8076 11200 8082 11212
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 8076 11172 9045 11200
rect 8076 11160 8082 11172
rect 9033 11169 9045 11172
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 9122 11160 9128 11212
rect 9180 11200 9186 11212
rect 9674 11200 9680 11212
rect 9180 11172 9680 11200
rect 9180 11160 9186 11172
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 9784 11172 12940 11200
rect 4338 11132 4344 11144
rect 4172 11104 4344 11132
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 7009 11135 7067 11141
rect 7009 11132 7021 11135
rect 5592 11104 7021 11132
rect 5592 11092 5598 11104
rect 7009 11101 7021 11104
rect 7055 11132 7067 11135
rect 7190 11132 7196 11144
rect 7055 11104 7196 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 7524 11104 7788 11132
rect 7524 11092 7530 11104
rect 2498 11024 2504 11076
rect 2556 11024 2562 11076
rect 4924 11067 4982 11073
rect 4924 11033 4936 11067
rect 4970 11064 4982 11067
rect 6086 11064 6092 11076
rect 4970 11036 6092 11064
rect 4970 11033 4982 11036
rect 4924 11027 4982 11033
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 6764 11067 6822 11073
rect 6764 11033 6776 11067
rect 6810 11064 6822 11067
rect 7650 11064 7656 11076
rect 6810 11036 7656 11064
rect 6810 11033 6822 11036
rect 6764 11027 6822 11033
rect 7650 11024 7656 11036
rect 7708 11024 7714 11076
rect 4706 10956 4712 11008
rect 4764 10996 4770 11008
rect 7466 10996 7472 11008
rect 4764 10968 7472 10996
rect 4764 10956 4770 10968
rect 7466 10956 7472 10968
rect 7524 10956 7530 11008
rect 7760 10996 7788 11104
rect 7834 11092 7840 11144
rect 7892 11092 7898 11144
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 9784 11132 9812 11172
rect 9640 11104 9812 11132
rect 9640 11092 9646 11104
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 10284 11104 10333 11132
rect 10284 11092 10290 11104
rect 10321 11101 10333 11104
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 10594 11092 10600 11144
rect 10652 11132 10658 11144
rect 10689 11135 10747 11141
rect 10689 11132 10701 11135
rect 10652 11104 10701 11132
rect 10652 11092 10658 11104
rect 10689 11101 10701 11104
rect 10735 11101 10747 11135
rect 11146 11132 11152 11144
rect 11107 11104 11152 11132
rect 10689 11095 10747 11101
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11101 11483 11135
rect 12250 11132 12256 11144
rect 12211 11104 12256 11132
rect 11425 11095 11483 11101
rect 7852 11064 7880 11092
rect 7852 11036 7972 11064
rect 7944 11005 7972 11036
rect 8386 11024 8392 11076
rect 8444 11064 8450 11076
rect 9309 11067 9367 11073
rect 9309 11064 9321 11067
rect 8444 11036 9321 11064
rect 8444 11024 8450 11036
rect 9309 11033 9321 11036
rect 9355 11033 9367 11067
rect 9309 11027 9367 11033
rect 10413 11067 10471 11073
rect 10413 11033 10425 11067
rect 10459 11033 10471 11067
rect 10413 11027 10471 11033
rect 10505 11067 10563 11073
rect 10505 11033 10517 11067
rect 10551 11064 10563 11067
rect 10778 11064 10784 11076
rect 10551 11036 10784 11064
rect 10551 11033 10563 11036
rect 10505 11027 10563 11033
rect 7837 10999 7895 11005
rect 7837 10996 7849 10999
rect 7760 10968 7849 10996
rect 7837 10965 7849 10968
rect 7883 10965 7895 10999
rect 7837 10959 7895 10965
rect 7929 10999 7987 11005
rect 7929 10965 7941 10999
rect 7975 10965 7987 10999
rect 7929 10959 7987 10965
rect 9217 10999 9275 11005
rect 9217 10965 9229 10999
rect 9263 10996 9275 10999
rect 9858 10996 9864 11008
rect 9263 10968 9864 10996
rect 9263 10965 9275 10968
rect 9217 10959 9275 10965
rect 9858 10956 9864 10968
rect 9916 10956 9922 11008
rect 10428 10996 10456 11027
rect 10778 11024 10784 11036
rect 10836 11024 10842 11076
rect 11440 11064 11468 11095
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 12710 11132 12716 11144
rect 12636 11104 12716 11132
rect 12526 11064 12532 11076
rect 11440 11036 12532 11064
rect 12526 11024 12532 11036
rect 12584 11064 12590 11076
rect 12636 11064 12664 11104
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12912 11141 12940 11172
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11101 12955 11135
rect 13538 11132 13544 11144
rect 13499 11104 13544 11132
rect 12897 11095 12955 11101
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 13354 11064 13360 11076
rect 12584 11036 12664 11064
rect 12728 11036 13360 11064
rect 12584 11024 12590 11036
rect 10870 10996 10876 11008
rect 10428 10968 10876 10996
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 11238 10996 11244 11008
rect 11199 10968 11244 10996
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 12066 10996 12072 11008
rect 12027 10968 12072 10996
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 12728 11005 12756 11036
rect 13354 11024 13360 11036
rect 13412 11024 13418 11076
rect 12713 10999 12771 11005
rect 12713 10965 12725 10999
rect 12759 10965 12771 10999
rect 12713 10959 12771 10965
rect 1104 10906 16836 10928
rect 1104 10854 4898 10906
rect 4950 10854 4962 10906
rect 5014 10854 5026 10906
rect 5078 10854 5090 10906
rect 5142 10854 5154 10906
rect 5206 10854 8846 10906
rect 8898 10854 8910 10906
rect 8962 10854 8974 10906
rect 9026 10854 9038 10906
rect 9090 10854 9102 10906
rect 9154 10854 12794 10906
rect 12846 10854 12858 10906
rect 12910 10854 12922 10906
rect 12974 10854 12986 10906
rect 13038 10854 13050 10906
rect 13102 10854 16836 10906
rect 1104 10832 16836 10854
rect 3510 10752 3516 10804
rect 3568 10792 3574 10804
rect 3605 10795 3663 10801
rect 3605 10792 3617 10795
rect 3568 10764 3617 10792
rect 3568 10752 3574 10764
rect 3605 10761 3617 10764
rect 3651 10761 3663 10795
rect 6546 10792 6552 10804
rect 3605 10755 3663 10761
rect 5460 10764 6552 10792
rect 4062 10724 4068 10736
rect 2898 10696 4068 10724
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 4246 10684 4252 10736
rect 4304 10724 4310 10736
rect 4718 10727 4776 10733
rect 4718 10724 4730 10727
rect 4304 10696 4730 10724
rect 4304 10684 4310 10696
rect 4718 10693 4730 10696
rect 4764 10724 4776 10727
rect 4890 10724 4896 10736
rect 4764 10696 4896 10724
rect 4764 10693 4776 10696
rect 4718 10687 4776 10693
rect 4890 10684 4896 10696
rect 4948 10684 4954 10736
rect 5460 10733 5488 10764
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 9585 10795 9643 10801
rect 8168 10764 9536 10792
rect 8168 10752 8174 10764
rect 5445 10727 5503 10733
rect 5445 10693 5457 10727
rect 5491 10693 5503 10727
rect 5445 10687 5503 10693
rect 5661 10727 5719 10733
rect 5661 10693 5673 10727
rect 5707 10724 5719 10727
rect 5902 10724 5908 10736
rect 5707 10696 5908 10724
rect 5707 10693 5719 10696
rect 5661 10687 5719 10693
rect 5902 10684 5908 10696
rect 5960 10684 5966 10736
rect 6362 10684 6368 10736
rect 6420 10724 6426 10736
rect 8472 10727 8530 10733
rect 6420 10696 8248 10724
rect 6420 10684 6426 10696
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 8220 10665 8248 10696
rect 8472 10693 8484 10727
rect 8518 10724 8530 10727
rect 9306 10724 9312 10736
rect 8518 10696 9312 10724
rect 8518 10693 8530 10696
rect 8472 10687 8530 10693
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 6621 10659 6679 10665
rect 6621 10656 6633 10659
rect 5408 10628 6633 10656
rect 5408 10616 5414 10628
rect 6621 10625 6633 10628
rect 6667 10625 6679 10659
rect 6621 10619 6679 10625
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8294 10616 8300 10668
rect 8352 10616 8358 10668
rect 9508 10656 9536 10764
rect 9585 10761 9597 10795
rect 9631 10792 9643 10795
rect 9674 10792 9680 10804
rect 9631 10764 9680 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 9824 10764 11529 10792
rect 9824 10752 9830 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 12158 10752 12164 10804
rect 12216 10792 12222 10804
rect 14090 10792 14096 10804
rect 12216 10764 14096 10792
rect 12216 10752 12222 10764
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 10778 10724 10784 10736
rect 10520 10696 10784 10724
rect 10318 10656 10324 10668
rect 9508 10628 10324 10656
rect 10318 10616 10324 10628
rect 10376 10616 10382 10668
rect 10413 10659 10471 10665
rect 10413 10652 10425 10659
rect 10459 10652 10471 10659
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10557 1455 10591
rect 1670 10588 1676 10600
rect 1631 10560 1676 10588
rect 1397 10551 1455 10557
rect 1412 10452 1440 10551
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 4985 10591 5043 10597
rect 4985 10557 4997 10591
rect 5031 10588 5043 10591
rect 5442 10588 5448 10600
rect 5031 10560 5448 10588
rect 5031 10557 5043 10560
rect 4985 10551 5043 10557
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 6362 10588 6368 10600
rect 6323 10560 6368 10588
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 8312 10588 8340 10616
rect 10410 10600 10416 10652
rect 10468 10600 10474 10652
rect 10226 10588 10232 10600
rect 7760 10560 8340 10588
rect 10187 10560 10232 10588
rect 3510 10520 3516 10532
rect 2746 10492 3516 10520
rect 2746 10452 2774 10492
rect 3510 10480 3516 10492
rect 3568 10480 3574 10532
rect 6270 10520 6276 10532
rect 5644 10492 6276 10520
rect 1412 10424 2774 10452
rect 3145 10455 3203 10461
rect 3145 10421 3157 10455
rect 3191 10452 3203 10455
rect 4246 10452 4252 10464
rect 3191 10424 4252 10452
rect 3191 10421 3203 10424
rect 3145 10415 3203 10421
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 5644 10461 5672 10492
rect 6270 10480 6276 10492
rect 6328 10480 6334 10532
rect 7466 10480 7472 10532
rect 7524 10520 7530 10532
rect 7760 10529 7788 10560
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 10520 10597 10548 10696
rect 10778 10684 10784 10696
rect 10836 10684 10842 10736
rect 11238 10684 11244 10736
rect 11296 10724 11302 10736
rect 12066 10724 12072 10736
rect 11296 10696 12072 10724
rect 11296 10684 11302 10696
rect 12066 10684 12072 10696
rect 12124 10684 12130 10736
rect 12342 10684 12348 10736
rect 12400 10724 12406 10736
rect 13906 10724 13912 10736
rect 12400 10696 13400 10724
rect 13867 10696 13912 10724
rect 12400 10684 12406 10696
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11440 10628 11713 10656
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10557 10563 10591
rect 10505 10551 10563 10557
rect 11440 10532 11468 10628
rect 11701 10625 11713 10628
rect 11747 10656 11759 10659
rect 12250 10656 12256 10668
rect 11747 10628 12256 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 12434 10656 12440 10668
rect 12395 10628 12440 10656
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10625 12587 10659
rect 12710 10656 12716 10668
rect 12671 10628 12716 10656
rect 12529 10619 12587 10625
rect 11977 10591 12035 10597
rect 11977 10588 11989 10591
rect 11532 10560 11989 10588
rect 7745 10523 7803 10529
rect 7745 10520 7757 10523
rect 7524 10492 7757 10520
rect 7524 10480 7530 10492
rect 7745 10489 7757 10492
rect 7791 10489 7803 10523
rect 7745 10483 7803 10489
rect 9876 10492 11376 10520
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10421 5687 10455
rect 5629 10415 5687 10421
rect 5813 10455 5871 10461
rect 5813 10421 5825 10455
rect 5859 10452 5871 10455
rect 9876 10452 9904 10492
rect 10042 10452 10048 10464
rect 5859 10424 9904 10452
rect 10003 10424 10048 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 11348 10452 11376 10492
rect 11422 10480 11428 10532
rect 11480 10480 11486 10532
rect 11532 10452 11560 10560
rect 11977 10557 11989 10560
rect 12023 10557 12035 10591
rect 11977 10551 12035 10557
rect 12066 10548 12072 10600
rect 12124 10588 12130 10600
rect 12544 10588 12572 10619
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 13170 10656 13176 10668
rect 13131 10628 13176 10656
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 13372 10665 13400 10696
rect 13906 10684 13912 10696
rect 13964 10684 13970 10736
rect 13357 10659 13415 10665
rect 13357 10625 13369 10659
rect 13403 10625 13415 10659
rect 13814 10656 13820 10668
rect 13775 10628 13820 10656
rect 13357 10619 13415 10625
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 14001 10659 14059 10665
rect 14001 10625 14013 10659
rect 14047 10625 14059 10659
rect 14642 10656 14648 10668
rect 14603 10628 14648 10656
rect 14001 10619 14059 10625
rect 12124 10560 12572 10588
rect 12124 10548 12130 10560
rect 13262 10548 13268 10600
rect 13320 10588 13326 10600
rect 14016 10588 14044 10619
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 13320 10560 14044 10588
rect 13320 10548 13326 10560
rect 11885 10523 11943 10529
rect 11885 10489 11897 10523
rect 11931 10520 11943 10523
rect 13173 10523 13231 10529
rect 13173 10520 13185 10523
rect 11931 10492 13185 10520
rect 11931 10489 11943 10492
rect 11885 10483 11943 10489
rect 13173 10489 13185 10492
rect 13219 10489 13231 10523
rect 13173 10483 13231 10489
rect 11348 10424 11560 10452
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 12710 10452 12716 10464
rect 12308 10424 12716 10452
rect 12308 10412 12314 10424
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 14458 10452 14464 10464
rect 14419 10424 14464 10452
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 1104 10362 16836 10384
rect 1104 10310 2924 10362
rect 2976 10310 2988 10362
rect 3040 10310 3052 10362
rect 3104 10310 3116 10362
rect 3168 10310 3180 10362
rect 3232 10310 6872 10362
rect 6924 10310 6936 10362
rect 6988 10310 7000 10362
rect 7052 10310 7064 10362
rect 7116 10310 7128 10362
rect 7180 10310 10820 10362
rect 10872 10310 10884 10362
rect 10936 10310 10948 10362
rect 11000 10310 11012 10362
rect 11064 10310 11076 10362
rect 11128 10310 14768 10362
rect 14820 10310 14832 10362
rect 14884 10310 14896 10362
rect 14948 10310 14960 10362
rect 15012 10310 15024 10362
rect 15076 10310 16836 10362
rect 1104 10288 16836 10310
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3752 10220 3801 10248
rect 3752 10208 3758 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 6362 10248 6368 10260
rect 3789 10211 3847 10217
rect 5644 10220 6368 10248
rect 5169 10115 5227 10121
rect 5169 10081 5181 10115
rect 5215 10112 5227 10115
rect 5534 10112 5540 10124
rect 5215 10084 5540 10112
rect 5215 10081 5227 10084
rect 5169 10075 5227 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 5644 10121 5672 10220
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 8113 10251 8171 10257
rect 8113 10248 8125 10251
rect 7340 10220 8125 10248
rect 7340 10208 7346 10220
rect 8113 10217 8125 10220
rect 8159 10217 8171 10251
rect 8113 10211 8171 10217
rect 10594 10208 10600 10260
rect 10652 10248 10658 10260
rect 10781 10251 10839 10257
rect 10781 10248 10793 10251
rect 10652 10220 10793 10248
rect 10652 10208 10658 10220
rect 10781 10217 10793 10220
rect 10827 10217 10839 10251
rect 10781 10211 10839 10217
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 11882 10248 11888 10260
rect 11572 10220 11888 10248
rect 11572 10208 11578 10220
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 14090 10248 14096 10260
rect 14051 10220 14096 10248
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 7009 10183 7067 10189
rect 7009 10149 7021 10183
rect 7055 10180 7067 10183
rect 8662 10180 8668 10192
rect 7055 10152 8668 10180
rect 7055 10149 7067 10152
rect 7009 10143 7067 10149
rect 8662 10140 8668 10152
rect 8720 10140 8726 10192
rect 9398 10140 9404 10192
rect 9456 10180 9462 10192
rect 11241 10183 11299 10189
rect 11241 10180 11253 10183
rect 9456 10152 11253 10180
rect 9456 10140 9462 10152
rect 11241 10149 11253 10152
rect 11287 10149 11299 10183
rect 11241 10143 11299 10149
rect 12250 10140 12256 10192
rect 12308 10180 12314 10192
rect 13173 10183 13231 10189
rect 13173 10180 13185 10183
rect 12308 10152 13185 10180
rect 12308 10140 12314 10152
rect 13173 10149 13185 10152
rect 13219 10149 13231 10183
rect 13173 10143 13231 10149
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 7834 10072 7840 10124
rect 7892 10112 7898 10124
rect 9033 10115 9091 10121
rect 9033 10112 9045 10115
rect 7892 10084 9045 10112
rect 7892 10072 7898 10084
rect 9033 10081 9045 10084
rect 9079 10081 9091 10115
rect 9033 10075 9091 10081
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 11517 10115 11575 10121
rect 11517 10112 11529 10115
rect 9548 10084 11529 10112
rect 9548 10072 9554 10084
rect 11517 10081 11529 10084
rect 11563 10081 11575 10115
rect 13262 10112 13268 10124
rect 11517 10075 11575 10081
rect 11624 10084 13268 10112
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10013 1547 10047
rect 1489 10007 1547 10013
rect 1504 9976 1532 10007
rect 4890 10004 4896 10056
rect 4948 10053 4954 10056
rect 4948 10044 4960 10053
rect 4948 10016 4993 10044
rect 4948 10007 4960 10016
rect 4948 10004 4954 10007
rect 6178 10004 6184 10056
rect 6236 10044 6242 10056
rect 7650 10053 7656 10056
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 6236 10016 7481 10044
rect 6236 10004 6242 10016
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7617 10047 7656 10053
rect 7617 10013 7629 10047
rect 7617 10007 7656 10013
rect 7650 10004 7656 10007
rect 7708 10004 7714 10056
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 7975 10047 8033 10053
rect 7800 10016 7845 10044
rect 7800 10004 7806 10016
rect 7975 10013 7987 10047
rect 8021 10044 8033 10047
rect 8294 10044 8300 10056
rect 8021 10016 8300 10044
rect 8021 10013 8033 10016
rect 7975 10007 8033 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9916 10016 10149 10044
rect 9916 10004 9922 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10137 10007 10195 10013
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10410 10004 10416 10056
rect 10468 10044 10474 10056
rect 10551 10047 10609 10053
rect 10468 10016 10513 10044
rect 10468 10004 10474 10016
rect 10551 10013 10563 10047
rect 10597 10044 10609 10047
rect 10778 10044 10784 10056
rect 10597 10016 10784 10044
rect 10597 10013 10609 10016
rect 10551 10007 10609 10013
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 11624 10053 11652 10084
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10013 11667 10047
rect 11609 10007 11667 10013
rect 1762 9976 1768 9988
rect 1504 9948 1624 9976
rect 1723 9948 1768 9976
rect 1596 9920 1624 9948
rect 1762 9936 1768 9948
rect 1820 9936 1826 9988
rect 3326 9976 3332 9988
rect 2990 9948 3332 9976
rect 3326 9936 3332 9948
rect 3384 9936 3390 9988
rect 4430 9976 4436 9988
rect 3528 9948 4436 9976
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 3237 9911 3295 9917
rect 3237 9877 3249 9911
rect 3283 9908 3295 9911
rect 3528 9908 3556 9948
rect 4430 9936 4436 9948
rect 4488 9936 4494 9988
rect 5874 9979 5932 9985
rect 5874 9976 5886 9979
rect 5000 9948 5886 9976
rect 3283 9880 3556 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 5000 9908 5028 9948
rect 5874 9945 5886 9948
rect 5920 9945 5932 9979
rect 5874 9939 5932 9945
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 7837 9979 7895 9985
rect 7837 9976 7849 9979
rect 6328 9948 7849 9976
rect 6328 9936 6334 9948
rect 7837 9945 7849 9948
rect 7883 9976 7895 9979
rect 9309 9979 9367 9985
rect 9309 9976 9321 9979
rect 7883 9948 9321 9976
rect 7883 9945 7895 9948
rect 7837 9939 7895 9945
rect 9309 9945 9321 9948
rect 9355 9976 9367 9979
rect 11624 9976 11652 10007
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 12253 10047 12311 10053
rect 12253 10044 12265 10047
rect 12124 10016 12265 10044
rect 12124 10004 12130 10016
rect 12253 10013 12265 10016
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10044 12587 10047
rect 12618 10044 12624 10056
rect 12575 10016 12624 10044
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 9355 9948 11652 9976
rect 9355 9945 9367 9948
rect 9309 9939 9367 9945
rect 3660 9880 5028 9908
rect 3660 9868 3666 9880
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 9217 9911 9275 9917
rect 9217 9908 9229 9911
rect 8444 9880 9229 9908
rect 8444 9868 8450 9880
rect 9217 9877 9229 9880
rect 9263 9877 9275 9911
rect 9217 9871 9275 9877
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 12360 9908 12388 10007
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 13357 10047 13415 10053
rect 13357 10044 13369 10047
rect 12768 10016 13369 10044
rect 12768 10004 12774 10016
rect 13357 10013 13369 10016
rect 13403 10013 13415 10047
rect 14274 10044 14280 10056
rect 14235 10016 14280 10044
rect 13357 10007 13415 10013
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 12710 9908 12716 9920
rect 9732 9880 12388 9908
rect 12671 9880 12716 9908
rect 9732 9868 9738 9880
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 1104 9818 16836 9840
rect 1104 9766 4898 9818
rect 4950 9766 4962 9818
rect 5014 9766 5026 9818
rect 5078 9766 5090 9818
rect 5142 9766 5154 9818
rect 5206 9766 8846 9818
rect 8898 9766 8910 9818
rect 8962 9766 8974 9818
rect 9026 9766 9038 9818
rect 9090 9766 9102 9818
rect 9154 9766 12794 9818
rect 12846 9766 12858 9818
rect 12910 9766 12922 9818
rect 12974 9766 12986 9818
rect 13038 9766 13050 9818
rect 13102 9766 16836 9818
rect 1104 9744 16836 9766
rect 1486 9664 1492 9716
rect 1544 9704 1550 9716
rect 1581 9707 1639 9713
rect 1581 9704 1593 9707
rect 1544 9676 1593 9704
rect 1544 9664 1550 9676
rect 1581 9673 1593 9676
rect 1627 9673 1639 9707
rect 1581 9667 1639 9673
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4304 9676 5304 9704
rect 4304 9664 4310 9676
rect 3970 9636 3976 9648
rect 2622 9608 3976 9636
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 5276 9645 5304 9676
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 5960 9676 7512 9704
rect 5960 9664 5966 9676
rect 5261 9639 5319 9645
rect 5261 9605 5273 9639
rect 5307 9636 5319 9639
rect 7374 9636 7380 9648
rect 5307 9608 7380 9636
rect 5307 9605 5319 9608
rect 5261 9599 5319 9605
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 7484 9636 7512 9676
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 9582 9704 9588 9716
rect 8168 9676 9588 9704
rect 8168 9664 8174 9676
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 9950 9704 9956 9716
rect 9695 9676 9956 9704
rect 9600 9636 9628 9664
rect 7484 9608 8340 9636
rect 4154 9528 4160 9580
rect 4212 9528 4218 9580
rect 6632 9571 6690 9577
rect 6632 9537 6644 9571
rect 6678 9568 6690 9571
rect 7190 9568 7196 9580
rect 6678 9540 7196 9568
rect 6678 9537 6690 9540
rect 6632 9531 6690 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3329 9503 3387 9509
rect 3099 9472 3280 9500
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3252 9432 3280 9472
rect 3329 9469 3341 9503
rect 3375 9500 3387 9503
rect 3694 9500 3700 9512
rect 3375 9472 3700 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 3694 9460 3700 9472
rect 3752 9460 3758 9512
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 5537 9503 5595 9509
rect 3844 9472 5488 9500
rect 3844 9460 3850 9472
rect 4246 9432 4252 9444
rect 3252 9404 4252 9432
rect 4246 9392 4252 9404
rect 4304 9392 4310 9444
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3476 9336 3801 9364
rect 3476 9324 3482 9336
rect 3789 9333 3801 9336
rect 3835 9364 3847 9367
rect 4798 9364 4804 9376
rect 3835 9336 4804 9364
rect 3835 9333 3847 9336
rect 3789 9327 3847 9333
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 5460 9364 5488 9472
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 6086 9500 6092 9512
rect 5583 9472 6092 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 6086 9460 6092 9472
rect 6144 9460 6150 9512
rect 6362 9500 6368 9512
rect 6323 9472 6368 9500
rect 6362 9460 6368 9472
rect 6420 9460 6426 9512
rect 7745 9435 7803 9441
rect 7745 9401 7757 9435
rect 7791 9432 7803 9435
rect 7926 9432 7932 9444
rect 7791 9404 7932 9432
rect 7791 9401 7803 9404
rect 7745 9395 7803 9401
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 8202 9432 8208 9444
rect 8163 9404 8208 9432
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 8312 9432 8340 9608
rect 9508 9608 9628 9636
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 8662 9568 8668 9580
rect 8527 9540 8668 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 9508 9577 9536 9608
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9568 8907 9571
rect 9493 9571 9551 9577
rect 8895 9540 9260 9568
rect 8895 9537 8907 9540
rect 8849 9531 8907 9537
rect 9232 9512 9260 9540
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9695 9558 9723 9676
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 12066 9704 12072 9716
rect 10284 9676 12072 9704
rect 10284 9664 10290 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 12434 9664 12440 9716
rect 12492 9664 12498 9716
rect 13265 9707 13323 9713
rect 13265 9673 13277 9707
rect 13311 9704 13323 9707
rect 13446 9704 13452 9716
rect 13311 9676 13452 9704
rect 13311 9673 13323 9676
rect 13265 9667 13323 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 9858 9636 9864 9648
rect 9819 9608 9864 9636
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 10597 9639 10655 9645
rect 10597 9605 10609 9639
rect 10643 9636 10655 9639
rect 11238 9636 11244 9648
rect 10643 9608 11244 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 12452 9636 12480 9664
rect 13354 9636 13360 9648
rect 11716 9608 12480 9636
rect 12636 9608 13360 9636
rect 10413 9571 10471 9577
rect 9968 9568 10180 9569
rect 10413 9568 10425 9571
rect 9600 9557 9723 9558
rect 9493 9531 9551 9537
rect 9585 9551 9723 9557
rect 9585 9517 9597 9551
rect 9631 9530 9723 9551
rect 9784 9541 10425 9568
rect 9784 9540 9996 9541
rect 10152 9540 10425 9541
rect 9631 9517 9643 9530
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8570 9500 8576 9512
rect 8435 9472 8576 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 8570 9460 8576 9472
rect 8628 9500 8634 9512
rect 9122 9500 9128 9512
rect 8628 9472 9128 9500
rect 8628 9460 8634 9472
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 9214 9460 9220 9512
rect 9272 9460 9278 9512
rect 9585 9511 9643 9517
rect 9784 9432 9812 9540
rect 10413 9537 10425 9540
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10502 9528 10508 9580
rect 10560 9568 10566 9580
rect 11716 9577 11744 9608
rect 12636 9580 12664 9608
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 10560 9540 10701 9568
rect 10560 9528 10566 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9537 11759 9571
rect 12342 9568 12348 9580
rect 12303 9540 12348 9568
rect 11701 9531 11759 9537
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9469 10011 9503
rect 9953 9463 10011 9469
rect 8312 9404 9812 9432
rect 9968 9432 9996 9463
rect 10594 9460 10600 9512
rect 10652 9500 10658 9512
rect 10796 9500 10824 9531
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12492 9540 12541 9568
rect 12492 9528 12498 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 13081 9571 13139 9577
rect 12676 9540 12721 9568
rect 12676 9528 12682 9540
rect 13081 9537 13093 9571
rect 13127 9537 13139 9571
rect 13262 9568 13268 9580
rect 13223 9540 13268 9568
rect 13081 9531 13139 9537
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 10652 9472 11529 9500
rect 10652 9460 10658 9472
rect 11517 9469 11529 9472
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11664 9472 11897 9500
rect 11664 9460 11670 9472
rect 11885 9469 11897 9472
rect 11931 9469 11943 9503
rect 13096 9500 13124 9531
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 11885 9463 11943 9469
rect 11992 9472 13124 9500
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 9968 9404 10977 9432
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 10965 9395 11023 9401
rect 11330 9392 11336 9444
rect 11388 9432 11394 9444
rect 11992 9432 12020 9472
rect 11388 9404 12020 9432
rect 11388 9392 11394 9404
rect 12066 9392 12072 9444
rect 12124 9432 12130 9444
rect 12437 9435 12495 9441
rect 12437 9432 12449 9435
rect 12124 9404 12449 9432
rect 12124 9392 12130 9404
rect 12437 9401 12449 9404
rect 12483 9401 12495 9435
rect 12437 9395 12495 9401
rect 6546 9364 6552 9376
rect 5460 9336 6552 9364
rect 6546 9324 6552 9336
rect 6604 9324 6610 9376
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 9309 9367 9367 9373
rect 9309 9364 9321 9367
rect 6696 9336 9321 9364
rect 6696 9324 6702 9336
rect 9309 9333 9321 9336
rect 9355 9333 9367 9367
rect 9309 9327 9367 9333
rect 9398 9324 9404 9376
rect 9456 9364 9462 9376
rect 14274 9364 14280 9376
rect 9456 9336 14280 9364
rect 9456 9324 9462 9336
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 1104 9274 16836 9296
rect 1104 9222 2924 9274
rect 2976 9222 2988 9274
rect 3040 9222 3052 9274
rect 3104 9222 3116 9274
rect 3168 9222 3180 9274
rect 3232 9222 6872 9274
rect 6924 9222 6936 9274
rect 6988 9222 7000 9274
rect 7052 9222 7064 9274
rect 7116 9222 7128 9274
rect 7180 9222 10820 9274
rect 10872 9222 10884 9274
rect 10936 9222 10948 9274
rect 11000 9222 11012 9274
rect 11064 9222 11076 9274
rect 11128 9222 14768 9274
rect 14820 9222 14832 9274
rect 14884 9222 14896 9274
rect 14948 9222 14960 9274
rect 15012 9222 15024 9274
rect 15076 9222 16836 9274
rect 1104 9200 16836 9222
rect 1443 9163 1501 9169
rect 1443 9129 1455 9163
rect 1489 9160 1501 9163
rect 1670 9160 1676 9172
rect 1489 9132 1676 9160
rect 1489 9129 1501 9132
rect 1443 9123 1501 9129
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 3016 9132 3924 9160
rect 3016 9120 3022 9132
rect 1578 8984 1584 9036
rect 1636 9024 1642 9036
rect 3789 9027 3847 9033
rect 3789 9024 3801 9027
rect 1636 8996 3801 9024
rect 1636 8984 1642 8996
rect 3789 8993 3801 8996
rect 3835 8993 3847 9027
rect 3896 9024 3924 9132
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 6454 9160 6460 9172
rect 4304 9132 6460 9160
rect 4304 9120 4310 9132
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 7837 9163 7895 9169
rect 7837 9160 7849 9163
rect 6604 9132 7849 9160
rect 6604 9120 6610 9132
rect 7837 9129 7849 9132
rect 7883 9129 7895 9163
rect 7837 9123 7895 9129
rect 7926 9120 7932 9172
rect 7984 9160 7990 9172
rect 9766 9160 9772 9172
rect 7984 9132 9772 9160
rect 7984 9120 7990 9132
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 10134 9160 10140 9172
rect 10095 9132 10140 9160
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10502 9120 10508 9172
rect 10560 9160 10566 9172
rect 10560 9132 11100 9160
rect 10560 9120 10566 9132
rect 5537 9095 5595 9101
rect 5537 9061 5549 9095
rect 5583 9092 5595 9095
rect 7282 9092 7288 9104
rect 5583 9064 7288 9092
rect 5583 9061 5595 9064
rect 5537 9055 5595 9061
rect 4522 9024 4528 9036
rect 3896 8996 4528 9024
rect 3789 8987 3847 8993
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 4614 8984 4620 9036
rect 4672 9024 4678 9036
rect 5552 9024 5580 9055
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 7650 9052 7656 9104
rect 7708 9092 7714 9104
rect 7745 9095 7803 9101
rect 7745 9092 7757 9095
rect 7708 9064 7757 9092
rect 7708 9052 7714 9064
rect 7745 9061 7757 9064
rect 7791 9061 7803 9095
rect 9582 9092 9588 9104
rect 7745 9055 7803 9061
rect 7852 9064 9588 9092
rect 6270 9024 6276 9036
rect 4672 8996 5580 9024
rect 6231 8996 6276 9024
rect 4672 8984 4678 8996
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 7852 9024 7880 9064
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 10594 9092 10600 9104
rect 10336 9064 10600 9092
rect 6380 8996 7880 9024
rect 7944 8996 8432 9024
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8956 2927 8959
rect 3237 8959 3295 8965
rect 2915 8928 3188 8956
rect 2915 8925 2927 8928
rect 2869 8919 2927 8925
rect 2314 8848 2320 8900
rect 2372 8848 2378 8900
rect 3160 8888 3188 8928
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 3510 8956 3516 8968
rect 3283 8928 3516 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 3418 8888 3424 8900
rect 3160 8860 3424 8888
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 4065 8891 4123 8897
rect 4065 8857 4077 8891
rect 4111 8857 4123 8891
rect 5442 8888 5448 8900
rect 5290 8860 5448 8888
rect 4065 8851 4123 8857
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 2958 8820 2964 8832
rect 1728 8792 2964 8820
rect 1728 8780 1734 8792
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 4080 8820 4108 8851
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 6012 8888 6040 8919
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 6380 8956 6408 8996
rect 6144 8928 6408 8956
rect 6144 8916 6150 8928
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7524 8928 7573 8956
rect 7524 8916 7530 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 7944 8956 7972 8996
rect 7699 8928 7972 8956
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 6270 8888 6276 8900
rect 6012 8860 6276 8888
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 5902 8820 5908 8832
rect 4080 8792 5908 8820
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 7285 8823 7343 8829
rect 7285 8789 7297 8823
rect 7331 8820 7343 8823
rect 7466 8820 7472 8832
rect 7331 8792 7472 8820
rect 7331 8789 7343 8792
rect 7285 8783 7343 8789
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 7576 8820 7604 8919
rect 7742 8820 7748 8832
rect 7576 8792 7748 8820
rect 7742 8780 7748 8792
rect 7800 8780 7806 8832
rect 7944 8820 7972 8928
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8956 8079 8959
rect 8202 8956 8208 8968
rect 8067 8928 8208 8956
rect 8067 8925 8079 8928
rect 8021 8919 8079 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8404 8956 8432 8996
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 8536 8996 9352 9024
rect 8536 8984 8542 8996
rect 8570 8956 8576 8968
rect 8404 8928 8576 8956
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 9122 8956 9128 8968
rect 9083 8928 9128 8956
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 9324 8965 9352 8996
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8925 9367 8959
rect 9490 8956 9496 8968
rect 9451 8928 9496 8956
rect 9309 8919 9367 8925
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9217 8891 9275 8897
rect 9217 8888 9229 8891
rect 9088 8860 9229 8888
rect 9088 8848 9094 8860
rect 9217 8857 9229 8860
rect 9263 8857 9275 8891
rect 10336 8888 10364 9064
rect 10594 9052 10600 9064
rect 10652 9052 10658 9104
rect 11072 9092 11100 9132
rect 11146 9120 11152 9172
rect 11204 9160 11210 9172
rect 12529 9163 12587 9169
rect 12529 9160 12541 9163
rect 11204 9132 12541 9160
rect 11204 9120 11210 9132
rect 12529 9129 12541 9132
rect 12575 9129 12587 9163
rect 12529 9123 12587 9129
rect 12618 9092 12624 9104
rect 11072 9064 12624 9092
rect 12618 9052 12624 9064
rect 12676 9052 12682 9104
rect 11054 8984 11060 9036
rect 11112 9024 11118 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 11112 8996 11161 9024
rect 11112 8984 11118 8996
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 12066 9024 12072 9036
rect 11149 8987 11207 8993
rect 11256 8996 12072 9024
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8956 10563 8959
rect 10594 8956 10600 8968
rect 10551 8928 10600 8956
rect 10551 8925 10563 8928
rect 10505 8919 10563 8925
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 11256 8956 11284 8996
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 10965 8919 11023 8925
rect 11072 8928 11284 8956
rect 9217 8851 9275 8857
rect 9324 8860 10364 8888
rect 9324 8832 9352 8860
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 10980 8888 11008 8919
rect 10468 8860 11008 8888
rect 10468 8848 10474 8860
rect 11072 8832 11100 8928
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 11974 8956 11980 8968
rect 11388 8928 11433 8956
rect 11935 8928 11980 8956
rect 11388 8916 11394 8928
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8925 12495 8959
rect 12618 8956 12624 8968
rect 12579 8928 12624 8956
rect 12437 8919 12495 8925
rect 11146 8848 11152 8900
rect 11204 8888 11210 8900
rect 12452 8888 12480 8919
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 11204 8860 12480 8888
rect 11204 8848 11210 8860
rect 8018 8820 8024 8832
rect 7944 8792 8024 8820
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8536 8792 8953 8820
rect 8536 8780 8542 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 9306 8780 9312 8832
rect 9364 8780 9370 8832
rect 9953 8823 10011 8829
rect 9953 8789 9965 8823
rect 9999 8820 10011 8823
rect 10042 8820 10048 8832
rect 9999 8792 10048 8820
rect 9999 8789 10011 8792
rect 9953 8783 10011 8789
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 10137 8823 10195 8829
rect 10137 8789 10149 8823
rect 10183 8820 10195 8823
rect 10502 8820 10508 8832
rect 10183 8792 10508 8820
rect 10183 8789 10195 8792
rect 10137 8783 10195 8789
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 11054 8820 11060 8832
rect 11015 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11238 8820 11244 8832
rect 11199 8792 11244 8820
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 11698 8780 11704 8832
rect 11756 8820 11762 8832
rect 11793 8823 11851 8829
rect 11793 8820 11805 8823
rect 11756 8792 11805 8820
rect 11756 8780 11762 8792
rect 11793 8789 11805 8792
rect 11839 8789 11851 8823
rect 11793 8783 11851 8789
rect 1104 8730 16836 8752
rect 1104 8678 4898 8730
rect 4950 8678 4962 8730
rect 5014 8678 5026 8730
rect 5078 8678 5090 8730
rect 5142 8678 5154 8730
rect 5206 8678 8846 8730
rect 8898 8678 8910 8730
rect 8962 8678 8974 8730
rect 9026 8678 9038 8730
rect 9090 8678 9102 8730
rect 9154 8678 12794 8730
rect 12846 8678 12858 8730
rect 12910 8678 12922 8730
rect 12974 8678 12986 8730
rect 13038 8678 13050 8730
rect 13102 8678 16836 8730
rect 1104 8656 16836 8678
rect 6822 8616 6828 8628
rect 3068 8588 6828 8616
rect 3068 8548 3096 8588
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7558 8616 7564 8628
rect 7147 8588 7564 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 9490 8616 9496 8628
rect 8036 8588 9496 8616
rect 2806 8520 3096 8548
rect 3191 8551 3249 8557
rect 3191 8517 3203 8551
rect 3237 8548 3249 8551
rect 3973 8551 4031 8557
rect 3973 8548 3985 8551
rect 3237 8520 3985 8548
rect 3237 8517 3249 8520
rect 3191 8511 3249 8517
rect 3973 8517 3985 8520
rect 4019 8517 4031 8551
rect 5258 8548 5264 8560
rect 5198 8520 5264 8548
rect 3973 8511 4031 8517
rect 5258 8508 5264 8520
rect 5316 8508 5322 8560
rect 8036 8548 8064 8588
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 9766 8616 9772 8628
rect 9727 8588 9772 8616
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 10502 8616 10508 8628
rect 10060 8588 10508 8616
rect 6656 8520 8064 8548
rect 8205 8551 8263 8557
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 6656 8489 6684 8520
rect 8205 8517 8217 8551
rect 8251 8548 8263 8551
rect 8478 8548 8484 8560
rect 8251 8520 8484 8548
rect 8251 8517 8263 8520
rect 8205 8511 8263 8517
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 9030 8508 9036 8560
rect 9088 8548 9094 8560
rect 10060 8548 10088 8588
rect 10502 8576 10508 8588
rect 10560 8616 10566 8628
rect 11701 8619 11759 8625
rect 11701 8616 11713 8619
rect 10560 8588 11713 8616
rect 10560 8576 10566 8588
rect 11701 8585 11713 8588
rect 11747 8616 11759 8619
rect 11790 8616 11796 8628
rect 11747 8588 11796 8616
rect 11747 8585 11759 8588
rect 11701 8579 11759 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 12158 8616 12164 8628
rect 12119 8588 12164 8616
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 10962 8548 10968 8560
rect 9088 8520 9260 8548
rect 9088 8508 9094 8520
rect 3697 8483 3755 8489
rect 3697 8480 3709 8483
rect 3568 8452 3709 8480
rect 3568 8440 3574 8452
rect 3697 8449 3709 8452
rect 3743 8449 3755 8483
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 3697 8443 3755 8449
rect 6380 8452 6653 8480
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8412 1823 8415
rect 1811 8384 3648 8412
rect 1811 8381 1823 8384
rect 1765 8375 1823 8381
rect 3620 8276 3648 8384
rect 4706 8372 4712 8424
rect 4764 8412 4770 8424
rect 6380 8412 6408 8452
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 6788 8452 6833 8480
rect 6788 8440 6794 8452
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7156 8452 7849 8480
rect 7156 8440 7162 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8662 8480 8668 8492
rect 8159 8452 8668 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 6546 8412 6552 8424
rect 4764 8384 6408 8412
rect 6472 8384 6552 8412
rect 4764 8372 4770 8384
rect 5074 8304 5080 8356
rect 5132 8344 5138 8356
rect 5445 8347 5503 8353
rect 5445 8344 5457 8347
rect 5132 8316 5457 8344
rect 5132 8304 5138 8316
rect 5445 8313 5457 8316
rect 5491 8313 5503 8347
rect 5445 8307 5503 8313
rect 5994 8304 6000 8356
rect 6052 8344 6058 8356
rect 6472 8344 6500 8384
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 8036 8412 8064 8440
rect 7791 8384 8064 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 7558 8344 7564 8356
rect 6052 8316 6500 8344
rect 7519 8316 7564 8344
rect 6052 8304 6058 8316
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 8018 8304 8024 8356
rect 8076 8344 8082 8356
rect 8128 8344 8156 8443
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8938 8480 8944 8492
rect 8899 8452 8944 8480
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 9232 8489 9260 8520
rect 9508 8520 10088 8548
rect 10336 8520 10548 8548
rect 9508 8492 9536 8520
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8480 9735 8483
rect 9766 8480 9772 8492
rect 9723 8452 9772 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 9933 8483 9991 8489
rect 9933 8449 9945 8483
rect 9979 8480 9991 8483
rect 10336 8480 10364 8520
rect 9979 8478 10088 8480
rect 10244 8478 10364 8480
rect 9979 8452 10364 8478
rect 9979 8450 9996 8452
rect 10060 8450 10272 8452
rect 9979 8449 9991 8450
rect 9933 8443 9991 8449
rect 10410 8412 10416 8424
rect 8076 8316 8156 8344
rect 8220 8384 10416 8412
rect 8076 8304 8082 8316
rect 4706 8276 4712 8288
rect 3620 8248 4712 8276
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 8220 8276 8248 8384
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 10520 8412 10548 8520
rect 10612 8520 10968 8548
rect 10612 8489 10640 8520
rect 10962 8508 10968 8520
rect 11020 8548 11026 8560
rect 11422 8548 11428 8560
rect 11020 8520 11428 8548
rect 11020 8508 11026 8520
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10686 8440 10692 8492
rect 10744 8478 10750 8492
rect 10781 8483 10839 8489
rect 10781 8478 10793 8483
rect 10744 8450 10793 8478
rect 10744 8440 10750 8450
rect 10781 8449 10793 8450
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 10928 8452 11529 8480
rect 10928 8440 10934 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 12161 8483 12219 8489
rect 12161 8480 12173 8483
rect 11664 8452 12173 8480
rect 11664 8440 11670 8452
rect 12161 8449 12173 8452
rect 12207 8449 12219 8483
rect 12342 8480 12348 8492
rect 12303 8452 12348 8480
rect 12161 8443 12219 8449
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 10965 8415 11023 8421
rect 10520 8384 10640 8412
rect 8662 8344 8668 8356
rect 8623 8316 8668 8344
rect 8662 8304 8668 8316
rect 8720 8304 8726 8356
rect 8754 8304 8760 8356
rect 8812 8344 8818 8356
rect 10137 8347 10195 8353
rect 8812 8316 9628 8344
rect 8812 8304 8818 8316
rect 6604 8248 8248 8276
rect 9125 8279 9183 8285
rect 6604 8236 6610 8248
rect 9125 8245 9137 8279
rect 9171 8276 9183 8279
rect 9490 8276 9496 8288
rect 9171 8248 9496 8276
rect 9171 8245 9183 8248
rect 9125 8239 9183 8245
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 9600 8276 9628 8316
rect 10137 8313 10149 8347
rect 10183 8344 10195 8347
rect 10502 8344 10508 8356
rect 10183 8316 10508 8344
rect 10183 8313 10195 8316
rect 10137 8307 10195 8313
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 10612 8344 10640 8384
rect 10965 8381 10977 8415
rect 11011 8412 11023 8415
rect 14642 8412 14648 8424
rect 11011 8384 14648 8412
rect 11011 8381 11023 8384
rect 10965 8375 11023 8381
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 12434 8344 12440 8356
rect 10612 8316 12440 8344
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 10778 8276 10784 8288
rect 9600 8248 10784 8276
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11238 8276 11244 8288
rect 11112 8248 11244 8276
rect 11112 8236 11118 8248
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 1104 8186 16836 8208
rect 1104 8134 2924 8186
rect 2976 8134 2988 8186
rect 3040 8134 3052 8186
rect 3104 8134 3116 8186
rect 3168 8134 3180 8186
rect 3232 8134 6872 8186
rect 6924 8134 6936 8186
rect 6988 8134 7000 8186
rect 7052 8134 7064 8186
rect 7116 8134 7128 8186
rect 7180 8134 10820 8186
rect 10872 8134 10884 8186
rect 10936 8134 10948 8186
rect 11000 8134 11012 8186
rect 11064 8134 11076 8186
rect 11128 8134 14768 8186
rect 14820 8134 14832 8186
rect 14884 8134 14896 8186
rect 14948 8134 14960 8186
rect 15012 8134 15024 8186
rect 15076 8134 16836 8186
rect 1104 8112 16836 8134
rect 3145 8075 3203 8081
rect 3145 8041 3157 8075
rect 3191 8072 3203 8075
rect 4246 8072 4252 8084
rect 3191 8044 4252 8072
rect 3191 8041 3203 8044
rect 3145 8035 3203 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4706 8032 4712 8084
rect 4764 8072 4770 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 4764 8044 5549 8072
rect 4764 8032 4770 8044
rect 5537 8041 5549 8044
rect 5583 8072 5595 8075
rect 7561 8075 7619 8081
rect 5583 8044 7521 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 6733 8007 6791 8013
rect 5920 7976 6500 8004
rect 3234 7896 3240 7948
rect 3292 7936 3298 7948
rect 5920 7936 5948 7976
rect 3292 7908 5948 7936
rect 3292 7896 3298 7908
rect 5994 7896 6000 7948
rect 6052 7936 6058 7948
rect 6181 7939 6239 7945
rect 6181 7936 6193 7939
rect 6052 7908 6193 7936
rect 6052 7896 6058 7908
rect 6181 7905 6193 7908
rect 6227 7905 6239 7939
rect 6181 7899 6239 7905
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1412 7732 1440 7831
rect 2774 7828 2780 7880
rect 2832 7828 2838 7880
rect 3786 7868 3792 7880
rect 3747 7840 3792 7868
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 6270 7868 6276 7880
rect 5684 7840 6276 7868
rect 5684 7828 5690 7840
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 6472 7868 6500 7976
rect 6733 7973 6745 8007
rect 6779 8004 6791 8007
rect 7098 8004 7104 8016
rect 6779 7976 7104 8004
rect 6779 7973 6791 7976
rect 6733 7967 6791 7973
rect 7098 7964 7104 7976
rect 7156 7964 7162 8016
rect 7493 8004 7521 8044
rect 7561 8041 7573 8075
rect 7607 8072 7619 8075
rect 7650 8072 7656 8084
rect 7607 8044 7656 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 7745 8075 7803 8081
rect 7745 8041 7757 8075
rect 7791 8072 7803 8075
rect 7834 8072 7840 8084
rect 7791 8044 7840 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 8294 8072 8300 8084
rect 8255 8044 8300 8072
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 10045 8075 10103 8081
rect 10045 8072 10057 8075
rect 9456 8044 10057 8072
rect 9456 8032 9462 8044
rect 10045 8041 10057 8044
rect 10091 8041 10103 8075
rect 11882 8072 11888 8084
rect 11843 8044 11888 8072
rect 10045 8035 10103 8041
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 8110 8004 8116 8016
rect 7493 7976 8116 8004
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 8478 7964 8484 8016
rect 8536 8004 8542 8016
rect 9033 8007 9091 8013
rect 9033 8004 9045 8007
rect 8536 7976 9045 8004
rect 8536 7964 8542 7976
rect 9033 7973 9045 7976
rect 9079 7973 9091 8007
rect 9033 7967 9091 7973
rect 9214 7964 9220 8016
rect 9272 8004 9278 8016
rect 13170 8004 13176 8016
rect 9272 7976 13176 8004
rect 9272 7964 9278 7976
rect 13170 7964 13176 7976
rect 13228 7964 13234 8016
rect 6822 7936 6828 7948
rect 6636 7908 6828 7936
rect 6636 7868 6664 7908
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 7892 7908 11253 7936
rect 7892 7896 7898 7908
rect 11241 7905 11253 7908
rect 11287 7905 11299 7939
rect 12434 7936 12440 7948
rect 11241 7899 11299 7905
rect 11348 7908 12440 7936
rect 6472 7840 6664 7868
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 7156 7840 7205 7868
rect 7156 7828 7162 7840
rect 7193 7837 7205 7840
rect 7239 7868 7251 7871
rect 7926 7868 7932 7880
rect 7239 7840 7932 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 8386 7868 8392 7880
rect 8299 7840 8392 7868
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 9858 7868 9864 7880
rect 9819 7840 9864 7868
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10502 7868 10508 7880
rect 10463 7840 10508 7868
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 10594 7828 10600 7880
rect 10652 7828 10658 7880
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7868 10747 7871
rect 10962 7868 10968 7880
rect 10735 7840 10968 7868
rect 10735 7837 10747 7840
rect 10689 7831 10747 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11146 7868 11152 7880
rect 11107 7840 11152 7868
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 11348 7877 11376 7908
rect 12434 7896 12440 7908
rect 12492 7936 12498 7948
rect 12618 7936 12624 7948
rect 12492 7908 12624 7936
rect 12492 7896 12498 7908
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11790 7868 11796 7880
rect 11751 7840 11796 7868
rect 11333 7831 11391 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 1670 7800 1676 7812
rect 1631 7772 1676 7800
rect 1670 7760 1676 7772
rect 1728 7760 1734 7812
rect 4062 7800 4068 7812
rect 4023 7772 4068 7800
rect 4062 7760 4068 7772
rect 4120 7760 4126 7812
rect 5442 7800 5448 7812
rect 5290 7772 5448 7800
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 6380 7800 6408 7828
rect 8404 7800 8432 7828
rect 9398 7800 9404 7812
rect 6380 7772 8432 7800
rect 9359 7772 9404 7800
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 10612 7800 10640 7828
rect 11992 7800 12020 7831
rect 10612 7772 12020 7800
rect 1578 7732 1584 7744
rect 1412 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 1688 7732 1716 7760
rect 2682 7732 2688 7744
rect 1688 7704 2688 7732
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 3510 7692 3516 7744
rect 3568 7732 3574 7744
rect 5074 7732 5080 7744
rect 3568 7704 5080 7732
rect 3568 7692 3574 7704
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6273 7735 6331 7741
rect 6273 7732 6285 7735
rect 5960 7704 6285 7732
rect 5960 7692 5966 7704
rect 6273 7701 6285 7704
rect 6319 7701 6331 7735
rect 6273 7695 6331 7701
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 7006 7732 7012 7744
rect 6420 7704 7012 7732
rect 6420 7692 6426 7704
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7340 7704 7573 7732
rect 7340 7692 7346 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8352 7704 8953 7732
rect 8352 7692 8358 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 8941 7695 8999 7701
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 10597 7735 10655 7741
rect 10597 7732 10609 7735
rect 9916 7704 10609 7732
rect 9916 7692 9922 7704
rect 10597 7701 10609 7704
rect 10643 7701 10655 7735
rect 10597 7695 10655 7701
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11238 7732 11244 7744
rect 11112 7704 11244 7732
rect 11112 7692 11118 7704
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 1104 7642 16836 7664
rect 1104 7590 4898 7642
rect 4950 7590 4962 7642
rect 5014 7590 5026 7642
rect 5078 7590 5090 7642
rect 5142 7590 5154 7642
rect 5206 7590 8846 7642
rect 8898 7590 8910 7642
rect 8962 7590 8974 7642
rect 9026 7590 9038 7642
rect 9090 7590 9102 7642
rect 9154 7590 12794 7642
rect 12846 7590 12858 7642
rect 12910 7590 12922 7642
rect 12974 7590 12986 7642
rect 13038 7590 13050 7642
rect 13102 7590 16836 7642
rect 1104 7568 16836 7590
rect 3510 7528 3516 7540
rect 1504 7500 3516 7528
rect 1504 7404 1532 7500
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 6917 7531 6975 7537
rect 3620 7500 6500 7528
rect 3234 7460 3240 7472
rect 2990 7432 3240 7460
rect 3234 7420 3240 7432
rect 3292 7420 3298 7472
rect 3620 7460 3648 7500
rect 3344 7432 3648 7460
rect 1486 7392 1492 7404
rect 1399 7364 1492 7392
rect 1486 7352 1492 7364
rect 1544 7352 1550 7404
rect 3050 7352 3056 7404
rect 3108 7392 3114 7404
rect 3344 7392 3372 7432
rect 3878 7420 3884 7472
rect 3936 7420 3942 7472
rect 3108 7364 3372 7392
rect 3108 7352 3114 7364
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 3896 7392 3924 7420
rect 3970 7401 3976 7404
rect 3568 7364 3924 7392
rect 3568 7352 3574 7364
rect 3964 7355 3976 7401
rect 4028 7392 4034 7404
rect 5537 7395 5595 7401
rect 4028 7364 4064 7392
rect 3970 7352 3976 7355
rect 4028 7352 4034 7364
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 1762 7324 1768 7336
rect 1723 7296 1768 7324
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 3697 7327 3755 7333
rect 3697 7324 3709 7327
rect 2464 7296 3709 7324
rect 2464 7284 2470 7296
rect 3697 7293 3709 7296
rect 3743 7293 3755 7327
rect 5552 7324 5580 7355
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 5816 7395 5874 7401
rect 5684 7364 5729 7392
rect 5684 7352 5690 7364
rect 5816 7361 5828 7395
rect 5862 7382 5874 7395
rect 5902 7382 5908 7404
rect 5862 7361 5908 7382
rect 5816 7355 5908 7361
rect 5828 7354 5908 7355
rect 5902 7352 5908 7354
rect 5960 7352 5966 7404
rect 6472 7402 6500 7500
rect 6652 7500 6776 7528
rect 6652 7469 6680 7500
rect 6641 7463 6699 7469
rect 6641 7429 6653 7463
rect 6687 7429 6699 7463
rect 6748 7460 6776 7500
rect 6917 7497 6929 7531
rect 6963 7528 6975 7531
rect 7190 7528 7196 7540
rect 6963 7500 7196 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 8754 7528 8760 7540
rect 7340 7500 8515 7528
rect 8715 7500 8760 7528
rect 7340 7488 7346 7500
rect 6748 7432 6960 7460
rect 6641 7423 6699 7429
rect 6472 7401 6592 7402
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6472 7395 6607 7401
rect 6472 7374 6561 7395
rect 6365 7355 6423 7361
rect 6549 7361 6561 7374
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 5718 7324 5724 7336
rect 5552 7296 5724 7324
rect 3697 7287 3755 7293
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 6380 7324 6408 7355
rect 6730 7352 6736 7404
rect 6788 7401 6794 7404
rect 6788 7395 6815 7401
rect 6803 7361 6815 7395
rect 6932 7392 6960 7432
rect 7006 7420 7012 7472
rect 7064 7460 7070 7472
rect 8386 7460 8392 7472
rect 7064 7432 8392 7460
rect 7064 7420 7070 7432
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 8487 7460 8515 7500
rect 8754 7488 8760 7500
rect 8812 7488 8818 7540
rect 10226 7528 10232 7540
rect 9232 7500 10232 7528
rect 8487 7432 8892 7460
rect 7282 7392 7288 7404
rect 6932 7364 7288 7392
rect 6788 7355 6815 7361
rect 6788 7352 6794 7355
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 7650 7392 7656 7404
rect 7607 7364 7656 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 8754 7392 8760 7404
rect 8619 7364 8760 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 8864 7392 8892 7432
rect 8938 7420 8944 7472
rect 8996 7460 9002 7472
rect 9232 7460 9260 7500
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 10410 7488 10416 7540
rect 10468 7528 10474 7540
rect 10505 7531 10563 7537
rect 10505 7528 10517 7531
rect 10468 7500 10517 7528
rect 10468 7488 10474 7500
rect 10505 7497 10517 7500
rect 10551 7497 10563 7531
rect 10505 7491 10563 7497
rect 9674 7460 9680 7472
rect 8996 7432 9260 7460
rect 8996 7420 9002 7432
rect 9232 7399 9260 7432
rect 9416 7432 9680 7460
rect 9416 7401 9444 7432
rect 9674 7420 9680 7432
rect 9732 7420 9738 7472
rect 11606 7460 11612 7472
rect 9876 7432 11612 7460
rect 9225 7393 9283 7399
rect 8864 7364 9076 7392
rect 6454 7324 6460 7336
rect 6380 7296 6460 7324
rect 6454 7284 6460 7296
rect 6512 7284 6518 7336
rect 7466 7324 7472 7336
rect 7427 7296 7472 7324
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7324 7987 7327
rect 8938 7324 8944 7336
rect 7975 7296 8944 7324
rect 7975 7293 7987 7296
rect 7929 7287 7987 7293
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 9048 7324 9076 7364
rect 9225 7359 9237 7393
rect 9271 7359 9283 7393
rect 9225 7353 9283 7359
rect 9411 7395 9469 7401
rect 9411 7361 9423 7395
rect 9457 7361 9469 7395
rect 9411 7355 9469 7361
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 9876 7401 9904 7432
rect 11606 7420 11612 7432
rect 11664 7420 11670 7472
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 9824 7364 9873 7392
rect 9824 7352 9830 7364
rect 9861 7361 9873 7364
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10502 7392 10508 7404
rect 10100 7364 10364 7392
rect 10463 7364 10508 7392
rect 10100 7352 10106 7364
rect 10336 7324 10364 7364
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 10689 7395 10747 7401
rect 10689 7392 10701 7395
rect 10652 7364 10701 7392
rect 10652 7352 10658 7364
rect 10689 7361 10701 7364
rect 10735 7361 10747 7395
rect 10689 7355 10747 7361
rect 12342 7324 12348 7336
rect 9048 7296 9260 7324
rect 10336 7296 12348 7324
rect 4706 7216 4712 7268
rect 4764 7256 4770 7268
rect 5077 7259 5135 7265
rect 5077 7256 5089 7259
rect 4764 7228 5089 7256
rect 4764 7216 4770 7228
rect 5077 7225 5089 7228
rect 5123 7225 5135 7259
rect 5077 7219 5135 7225
rect 5813 7259 5871 7265
rect 5813 7225 5825 7259
rect 5859 7256 5871 7259
rect 9122 7256 9128 7268
rect 5859 7228 9128 7256
rect 5859 7225 5871 7228
rect 5813 7219 5871 7225
rect 9122 7216 9128 7228
rect 9180 7216 9186 7268
rect 9232 7256 9260 7296
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 12250 7256 12256 7268
rect 9232 7228 12256 7256
rect 12250 7216 12256 7228
rect 12308 7216 12314 7268
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 3050 7188 3056 7200
rect 2188 7160 3056 7188
rect 2188 7148 2194 7160
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 3237 7191 3295 7197
rect 3237 7157 3249 7191
rect 3283 7188 3295 7191
rect 3510 7188 3516 7200
rect 3283 7160 3516 7188
rect 3283 7157 3295 7160
rect 3237 7151 3295 7157
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 9309 7191 9367 7197
rect 9309 7188 9321 7191
rect 5040 7160 9321 7188
rect 5040 7148 5046 7160
rect 9309 7157 9321 7160
rect 9355 7157 9367 7191
rect 9309 7151 9367 7157
rect 9398 7148 9404 7200
rect 9456 7188 9462 7200
rect 9953 7191 10011 7197
rect 9953 7188 9965 7191
rect 9456 7160 9965 7188
rect 9456 7148 9462 7160
rect 9953 7157 9965 7160
rect 9999 7157 10011 7191
rect 9953 7151 10011 7157
rect 1104 7098 16836 7120
rect 1104 7046 2924 7098
rect 2976 7046 2988 7098
rect 3040 7046 3052 7098
rect 3104 7046 3116 7098
rect 3168 7046 3180 7098
rect 3232 7046 6872 7098
rect 6924 7046 6936 7098
rect 6988 7046 7000 7098
rect 7052 7046 7064 7098
rect 7116 7046 7128 7098
rect 7180 7046 10820 7098
rect 10872 7046 10884 7098
rect 10936 7046 10948 7098
rect 11000 7046 11012 7098
rect 11064 7046 11076 7098
rect 11128 7046 14768 7098
rect 14820 7046 14832 7098
rect 14884 7046 14896 7098
rect 14948 7046 14960 7098
rect 15012 7046 15024 7098
rect 15076 7046 16836 7098
rect 1104 7024 16836 7046
rect 1486 6944 1492 6996
rect 1544 6984 1550 6996
rect 1654 6987 1712 6993
rect 1654 6984 1666 6987
rect 1544 6956 1666 6984
rect 1544 6944 1550 6956
rect 1654 6953 1666 6956
rect 1700 6953 1712 6987
rect 1654 6947 1712 6953
rect 3145 6987 3203 6993
rect 3145 6953 3157 6987
rect 3191 6984 3203 6987
rect 4062 6984 4068 6996
rect 3191 6956 4068 6984
rect 3191 6953 3203 6956
rect 3145 6947 3203 6953
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 5166 6984 5172 6996
rect 5127 6956 5172 6984
rect 5166 6944 5172 6956
rect 5224 6944 5230 6996
rect 5626 6984 5632 6996
rect 5587 6956 5632 6984
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 5994 6984 6000 6996
rect 5736 6956 6000 6984
rect 2866 6876 2872 6928
rect 2924 6916 2930 6928
rect 3878 6916 3884 6928
rect 2924 6888 3884 6916
rect 2924 6876 2930 6888
rect 3878 6876 3884 6888
rect 3936 6876 3942 6928
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 5184 6916 5212 6944
rect 4212 6888 5212 6916
rect 4212 6876 4218 6888
rect 5534 6876 5540 6928
rect 5592 6916 5598 6928
rect 5736 6916 5764 6956
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 6086 6944 6092 6996
rect 6144 6984 6150 6996
rect 6144 6956 6189 6984
rect 6144 6944 6150 6956
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 6822 6984 6828 6996
rect 6420 6956 6828 6984
rect 6420 6944 6426 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 8754 6984 8760 6996
rect 7064 6956 8760 6984
rect 7064 6944 7070 6956
rect 8754 6944 8760 6956
rect 8812 6944 8818 6996
rect 9030 6984 9036 6996
rect 8991 6956 9036 6984
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 9582 6984 9588 6996
rect 9543 6956 9588 6984
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 5592 6888 5764 6916
rect 5592 6876 5598 6888
rect 6730 6876 6736 6928
rect 6788 6916 6794 6928
rect 9306 6916 9312 6928
rect 6788 6888 9312 6916
rect 6788 6876 6794 6888
rect 9306 6876 9312 6888
rect 9364 6876 9370 6928
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 3142 6808 3148 6860
rect 3200 6848 3206 6860
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 3200 6820 3801 6848
rect 3200 6808 3206 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 4062 6848 4068 6860
rect 4023 6820 4068 6848
rect 3789 6811 3847 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4430 6808 4436 6860
rect 4488 6848 4494 6860
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 4488 6820 5365 6848
rect 4488 6808 4494 6820
rect 5353 6817 5365 6820
rect 5399 6848 5411 6851
rect 6273 6851 6331 6857
rect 6273 6848 6285 6851
rect 5399 6820 6285 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 6273 6817 6285 6820
rect 6319 6848 6331 6851
rect 7466 6848 7472 6860
rect 6319 6820 7472 6848
rect 6319 6817 6331 6820
rect 6273 6811 6331 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 8662 6848 8668 6860
rect 7616 6820 7661 6848
rect 8220 6820 8668 6848
rect 7616 6808 7622 6820
rect 1412 6644 1440 6808
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4304 6752 5089 6780
rect 4304 6740 4310 6752
rect 5077 6749 5089 6752
rect 5123 6780 5135 6783
rect 6089 6783 6147 6789
rect 6089 6780 6101 6783
rect 5123 6752 6101 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 6089 6749 6101 6752
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6780 6423 6783
rect 6546 6780 6552 6792
rect 6411 6752 6552 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6972 6752 7113 6780
rect 6972 6740 6978 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 7742 6780 7748 6792
rect 7423 6752 7748 6780
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 7463 6746 7512 6752
rect 2898 6684 5212 6712
rect 3786 6644 3792 6656
rect 1412 6616 3792 6644
rect 3786 6604 3792 6616
rect 3844 6644 3850 6656
rect 4062 6644 4068 6656
rect 3844 6616 4068 6644
rect 3844 6604 3850 6616
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 4430 6604 4436 6656
rect 4488 6644 4494 6656
rect 4982 6644 4988 6656
rect 4488 6616 4988 6644
rect 4488 6604 4494 6616
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 5184 6644 5212 6684
rect 5810 6672 5816 6724
rect 5868 6712 5874 6724
rect 6730 6712 6736 6724
rect 5868 6684 6736 6712
rect 5868 6672 5874 6684
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 7006 6672 7012 6724
rect 7064 6712 7070 6724
rect 7208 6712 7236 6743
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 8220 6789 8248 6820
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 10134 6848 10140 6860
rect 9048 6820 10140 6848
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7984 6752 8033 6780
rect 7984 6740 7990 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 7064 6684 7236 6712
rect 7064 6672 7070 6684
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 8312 6712 8340 6743
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 8941 6783 8999 6789
rect 8444 6774 8708 6780
rect 8941 6774 8953 6783
rect 8444 6752 8953 6774
rect 8444 6740 8450 6752
rect 8680 6749 8953 6752
rect 8987 6749 8999 6783
rect 8680 6746 8999 6749
rect 8941 6743 8999 6746
rect 9048 6712 9076 6820
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6774 9183 6783
rect 9214 6774 9220 6792
rect 9171 6749 9220 6774
rect 9125 6746 9220 6749
rect 9125 6743 9183 6746
rect 9214 6740 9220 6746
rect 9272 6740 9278 6792
rect 9582 6780 9588 6792
rect 9543 6752 9588 6780
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6780 9830 6792
rect 11422 6780 11428 6792
rect 9824 6752 11428 6780
rect 9824 6740 9830 6752
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 8168 6684 9076 6712
rect 8168 6672 8174 6684
rect 5994 6644 6000 6656
rect 5184 6616 6000 6644
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 6270 6604 6276 6656
rect 6328 6644 6334 6656
rect 6454 6644 6460 6656
rect 6328 6616 6460 6644
rect 6328 6604 6334 6616
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 9950 6644 9956 6656
rect 6595 6616 9956 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 1104 6554 16836 6576
rect 1104 6502 4898 6554
rect 4950 6502 4962 6554
rect 5014 6502 5026 6554
rect 5078 6502 5090 6554
rect 5142 6502 5154 6554
rect 5206 6502 8846 6554
rect 8898 6502 8910 6554
rect 8962 6502 8974 6554
rect 9026 6502 9038 6554
rect 9090 6502 9102 6554
rect 9154 6502 12794 6554
rect 12846 6502 12858 6554
rect 12910 6502 12922 6554
rect 12974 6502 12986 6554
rect 13038 6502 13050 6554
rect 13102 6502 16836 6554
rect 1104 6480 16836 6502
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 4982 6440 4988 6452
rect 2832 6412 2877 6440
rect 4356 6412 4988 6440
rect 2832 6400 2838 6412
rect 1664 6375 1722 6381
rect 1664 6341 1676 6375
rect 1710 6372 1722 6375
rect 1854 6372 1860 6384
rect 1710 6344 1860 6372
rect 1710 6341 1722 6344
rect 1664 6335 1722 6341
rect 1854 6332 1860 6344
rect 1912 6332 1918 6384
rect 2406 6332 2412 6384
rect 2464 6372 2470 6384
rect 4356 6372 4384 6412
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 5077 6443 5135 6449
rect 5077 6409 5089 6443
rect 5123 6440 5135 6443
rect 5350 6440 5356 6452
rect 5123 6412 5356 6440
rect 5123 6409 5135 6412
rect 5077 6403 5135 6409
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 5721 6443 5779 6449
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 5810 6440 5816 6452
rect 5767 6412 5816 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 6362 6440 6368 6452
rect 6323 6412 6368 6440
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 7285 6443 7343 6449
rect 7285 6440 7297 6443
rect 6880 6412 7297 6440
rect 6880 6400 6886 6412
rect 7285 6409 7297 6412
rect 7331 6409 7343 6443
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 7285 6403 7343 6409
rect 7668 6412 8309 6440
rect 2464 6344 4384 6372
rect 2464 6332 2470 6344
rect 4430 6332 4436 6384
rect 4488 6372 4494 6384
rect 4706 6372 4712 6384
rect 4488 6344 4568 6372
rect 4667 6344 4712 6372
rect 4488 6332 4494 6344
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 1486 6304 1492 6316
rect 1443 6276 1492 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 1486 6264 1492 6276
rect 1544 6264 1550 6316
rect 1946 6264 1952 6316
rect 2004 6304 2010 6316
rect 3142 6304 3148 6316
rect 2004 6276 3148 6304
rect 2004 6264 2010 6276
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6304 3847 6307
rect 4246 6304 4252 6316
rect 3835 6276 4252 6304
rect 3835 6273 3847 6276
rect 3789 6267 3847 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4540 6313 4568 6344
rect 4706 6332 4712 6344
rect 4764 6332 4770 6384
rect 4801 6375 4859 6381
rect 4801 6341 4813 6375
rect 4847 6372 4859 6375
rect 5537 6375 5595 6381
rect 5537 6372 5549 6375
rect 4847 6344 5549 6372
rect 4847 6341 4859 6344
rect 4801 6335 4859 6341
rect 5537 6341 5549 6344
rect 5583 6341 5595 6375
rect 6086 6372 6092 6384
rect 5537 6335 5595 6341
rect 5736 6344 6092 6372
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 3160 6168 3188 6264
rect 3510 6196 3516 6248
rect 3568 6236 3574 6248
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 3568 6208 4077 6236
rect 3568 6196 3574 6208
rect 4065 6205 4077 6208
rect 4111 6236 4123 6239
rect 4338 6236 4344 6248
rect 4111 6208 4344 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 3786 6168 3792 6180
rect 3160 6140 3792 6168
rect 3786 6128 3792 6140
rect 3844 6128 3850 6180
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 4816 6100 4844 6335
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 4908 6236 4936 6267
rect 5074 6264 5080 6316
rect 5132 6264 5138 6316
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5626 6304 5632 6316
rect 5408 6276 5632 6304
rect 5408 6264 5414 6276
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 5736 6304 5764 6344
rect 6086 6332 6092 6344
rect 6144 6332 6150 6384
rect 6270 6332 6276 6384
rect 6328 6372 6334 6384
rect 7668 6381 7696 6412
rect 8297 6409 8309 6412
rect 8343 6440 8355 6443
rect 10686 6440 10692 6452
rect 8343 6412 10692 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 7437 6375 7495 6381
rect 7437 6372 7449 6375
rect 6328 6344 7449 6372
rect 6328 6332 6334 6344
rect 7437 6341 7449 6344
rect 7483 6341 7495 6375
rect 7437 6335 7495 6341
rect 7653 6375 7711 6381
rect 7653 6341 7665 6375
rect 7699 6341 7711 6375
rect 7653 6335 7711 6341
rect 5797 6307 5855 6313
rect 5797 6304 5809 6307
rect 5736 6276 5809 6304
rect 5797 6273 5809 6276
rect 5843 6273 5855 6307
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 5797 6267 5855 6273
rect 6012 6276 6561 6304
rect 4982 6236 4988 6248
rect 4908 6208 4988 6236
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5092 6236 5120 6264
rect 6012 6236 6040 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6304 6883 6307
rect 7190 6304 7196 6316
rect 6871 6276 7196 6304
rect 6871 6273 6883 6276
rect 6825 6267 6883 6273
rect 5092 6208 6040 6236
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 6748 6236 6776 6267
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 7300 6304 7420 6308
rect 7668 6304 7696 6335
rect 7742 6332 7748 6384
rect 7800 6372 7806 6384
rect 9214 6372 9220 6384
rect 7800 6344 9220 6372
rect 7800 6332 7806 6344
rect 9214 6332 9220 6344
rect 9272 6372 9278 6384
rect 10042 6372 10048 6384
rect 9272 6344 10048 6372
rect 9272 6332 9278 6344
rect 10042 6332 10048 6344
rect 10100 6332 10106 6384
rect 8110 6304 8116 6316
rect 7300 6280 7696 6304
rect 7300 6236 7328 6280
rect 7392 6276 7696 6280
rect 8071 6276 8116 6304
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8628 6276 8953 6304
rect 8628 6264 8634 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 6144 6208 7328 6236
rect 6144 6196 6150 6208
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 9582 6236 9588 6248
rect 8720 6208 9588 6236
rect 8720 6196 8726 6208
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 5074 6128 5080 6180
rect 5132 6168 5138 6180
rect 5537 6171 5595 6177
rect 5537 6168 5549 6171
rect 5132 6140 5549 6168
rect 5132 6128 5138 6140
rect 5537 6137 5549 6140
rect 5583 6137 5595 6171
rect 5537 6131 5595 6137
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 7834 6168 7840 6180
rect 6052 6140 7840 6168
rect 6052 6128 6058 6140
rect 7834 6128 7840 6140
rect 7892 6128 7898 6180
rect 8754 6168 8760 6180
rect 8715 6140 8760 6168
rect 8754 6128 8760 6140
rect 8812 6128 8818 6180
rect 7190 6100 7196 6112
rect 3568 6072 7196 6100
rect 3568 6060 3574 6072
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 7475 6060 7481 6112
rect 7533 6100 7539 6112
rect 7533 6072 7578 6100
rect 7533 6060 7539 6072
rect 8110 6060 8116 6112
rect 8168 6100 8174 6112
rect 11146 6100 11152 6112
rect 8168 6072 11152 6100
rect 8168 6060 8174 6072
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 1104 6010 16836 6032
rect 1104 5958 2924 6010
rect 2976 5958 2988 6010
rect 3040 5958 3052 6010
rect 3104 5958 3116 6010
rect 3168 5958 3180 6010
rect 3232 5958 6872 6010
rect 6924 5958 6936 6010
rect 6988 5958 7000 6010
rect 7052 5958 7064 6010
rect 7116 5958 7128 6010
rect 7180 5958 10820 6010
rect 10872 5958 10884 6010
rect 10936 5958 10948 6010
rect 11000 5958 11012 6010
rect 11064 5958 11076 6010
rect 11128 5958 14768 6010
rect 14820 5958 14832 6010
rect 14884 5958 14896 6010
rect 14948 5958 14960 6010
rect 15012 5958 15024 6010
rect 15076 5958 16836 6010
rect 1104 5936 16836 5958
rect 4522 5856 4528 5908
rect 4580 5896 4586 5908
rect 6273 5899 6331 5905
rect 6273 5896 6285 5899
rect 4580 5868 6285 5896
rect 4580 5856 4586 5868
rect 6273 5865 6285 5868
rect 6319 5865 6331 5899
rect 6273 5859 6331 5865
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 7653 5899 7711 5905
rect 7653 5896 7665 5899
rect 6604 5868 7665 5896
rect 6604 5856 6610 5868
rect 7653 5865 7665 5868
rect 7699 5865 7711 5899
rect 7653 5859 7711 5865
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 7558 5828 7564 5840
rect 3844 5800 7564 5828
rect 3844 5788 3850 5800
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 1762 5720 1768 5772
rect 1820 5760 1826 5772
rect 4065 5763 4123 5769
rect 1820 5732 3924 5760
rect 1820 5720 1826 5732
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5661 2467 5695
rect 2409 5655 2467 5661
rect 2424 5624 2452 5655
rect 2590 5652 2596 5704
rect 2648 5692 2654 5704
rect 2685 5695 2743 5701
rect 2685 5692 2697 5695
rect 2648 5664 2697 5692
rect 2648 5652 2654 5664
rect 2685 5661 2697 5664
rect 2731 5661 2743 5695
rect 3786 5692 3792 5704
rect 3747 5664 3792 5692
rect 2685 5655 2743 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 3896 5692 3924 5732
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 4522 5760 4528 5772
rect 4111 5732 4528 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 5169 5763 5227 5769
rect 5169 5760 5181 5763
rect 4816 5732 5181 5760
rect 4816 5692 4844 5732
rect 5169 5729 5181 5732
rect 5215 5760 5227 5763
rect 5626 5760 5632 5772
rect 5215 5732 5488 5760
rect 5587 5732 5632 5760
rect 5215 5729 5227 5732
rect 5169 5723 5227 5729
rect 5261 5695 5319 5701
rect 5261 5692 5273 5695
rect 3896 5664 4844 5692
rect 5184 5664 5273 5692
rect 3970 5624 3976 5636
rect 2424 5596 3976 5624
rect 3970 5584 3976 5596
rect 4028 5584 4034 5636
rect 4246 5584 4252 5636
rect 4304 5624 4310 5636
rect 5184 5624 5212 5664
rect 5261 5661 5273 5664
rect 5307 5692 5319 5695
rect 5350 5692 5356 5704
rect 5307 5664 5356 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5460 5692 5488 5732
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5760 7067 5763
rect 7282 5760 7288 5772
rect 7055 5732 7288 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 8478 5760 8484 5772
rect 7576 5732 8484 5760
rect 6730 5692 6736 5704
rect 5460 5664 6736 5692
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 6914 5692 6920 5704
rect 6875 5664 6920 5692
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 7374 5692 7380 5704
rect 7147 5664 7380 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 7374 5652 7380 5664
rect 7432 5652 7438 5704
rect 7576 5701 7604 5732
rect 8478 5720 8484 5732
rect 8536 5760 8542 5772
rect 9674 5760 9680 5772
rect 8536 5732 9680 5760
rect 8536 5720 8542 5732
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5661 7619 5695
rect 7742 5692 7748 5704
rect 7703 5664 7748 5692
rect 7561 5655 7619 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 7892 5664 8401 5692
rect 7892 5652 7898 5664
rect 8389 5661 8401 5664
rect 8435 5692 8447 5695
rect 10502 5692 10508 5704
rect 8435 5664 10508 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 6086 5624 6092 5636
rect 4304 5596 5212 5624
rect 6047 5596 6092 5624
rect 4304 5584 4310 5596
rect 6086 5584 6092 5596
rect 6144 5584 6150 5636
rect 10594 5624 10600 5636
rect 6196 5596 10600 5624
rect 2590 5516 2596 5568
rect 2648 5556 2654 5568
rect 6196 5556 6224 5596
rect 10594 5584 10600 5596
rect 10652 5584 10658 5636
rect 2648 5528 6224 5556
rect 2648 5516 2654 5528
rect 6270 5516 6276 5568
rect 6328 5565 6334 5568
rect 6328 5559 6347 5565
rect 6335 5525 6347 5559
rect 6328 5519 6347 5525
rect 6457 5559 6515 5565
rect 6457 5525 6469 5559
rect 6503 5556 6515 5559
rect 7098 5556 7104 5568
rect 6503 5528 7104 5556
rect 6503 5525 6515 5528
rect 6457 5519 6515 5525
rect 6328 5516 6334 5519
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7374 5516 7380 5568
rect 7432 5556 7438 5568
rect 8018 5556 8024 5568
rect 7432 5528 8024 5556
rect 7432 5516 7438 5528
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 8205 5559 8263 5565
rect 8205 5525 8217 5559
rect 8251 5556 8263 5559
rect 8478 5556 8484 5568
rect 8251 5528 8484 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 1104 5466 16836 5488
rect 1104 5414 4898 5466
rect 4950 5414 4962 5466
rect 5014 5414 5026 5466
rect 5078 5414 5090 5466
rect 5142 5414 5154 5466
rect 5206 5414 8846 5466
rect 8898 5414 8910 5466
rect 8962 5414 8974 5466
rect 9026 5414 9038 5466
rect 9090 5414 9102 5466
rect 9154 5414 12794 5466
rect 12846 5414 12858 5466
rect 12910 5414 12922 5466
rect 12974 5414 12986 5466
rect 13038 5414 13050 5466
rect 13102 5414 16836 5466
rect 1104 5392 16836 5414
rect 3602 5352 3608 5364
rect 3563 5324 3608 5352
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 5077 5355 5135 5361
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5350 5352 5356 5364
rect 5123 5324 5356 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 6270 5352 6276 5364
rect 5592 5324 6276 5352
rect 5592 5312 5598 5324
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 6454 5352 6460 5364
rect 6415 5324 6460 5352
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 7190 5352 7196 5364
rect 6972 5324 7196 5352
rect 6972 5312 6978 5324
rect 7190 5312 7196 5324
rect 7248 5352 7254 5364
rect 11974 5352 11980 5364
rect 7248 5324 11980 5352
rect 7248 5312 7254 5324
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 3329 5287 3387 5293
rect 3329 5253 3341 5287
rect 3375 5284 3387 5287
rect 3510 5284 3516 5296
rect 3375 5256 3516 5284
rect 3375 5253 3387 5256
rect 3329 5247 3387 5253
rect 3510 5244 3516 5256
rect 3568 5244 3574 5296
rect 5445 5287 5503 5293
rect 5215 5253 5273 5259
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5216 2375 5219
rect 2498 5216 2504 5228
rect 2363 5188 2504 5216
rect 2363 5185 2375 5188
rect 2317 5179 2375 5185
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 3050 5216 3056 5228
rect 3011 5188 3056 5216
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 3234 5216 3240 5228
rect 3195 5188 3240 5216
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5216 3479 5219
rect 3970 5216 3976 5228
rect 3467 5188 3976 5216
rect 3467 5185 3479 5188
rect 3421 5179 3479 5185
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4246 5216 4252 5228
rect 4207 5188 4252 5216
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 5215 5219 5227 5253
rect 5261 5250 5273 5253
rect 5445 5253 5457 5287
rect 5491 5284 5503 5287
rect 6086 5284 6092 5296
rect 5491 5256 6092 5284
rect 5491 5253 5503 5256
rect 5261 5219 5288 5250
rect 5445 5247 5503 5253
rect 6086 5244 6092 5256
rect 6144 5244 6150 5296
rect 8478 5284 8484 5296
rect 6564 5256 8484 5284
rect 5215 5216 5288 5219
rect 5534 5216 5540 5228
rect 5215 5213 5540 5216
rect 5260 5188 5540 5213
rect 5534 5176 5540 5188
rect 5592 5176 5598 5228
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 5776 5188 6040 5216
rect 5776 5176 5782 5188
rect 6012 5160 6040 5188
rect 6362 5176 6368 5228
rect 6420 5216 6426 5228
rect 6564 5225 6592 5256
rect 8478 5244 8484 5256
rect 8536 5244 8542 5296
rect 6549 5219 6607 5225
rect 6420 5188 6465 5216
rect 6420 5176 6426 5188
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 6788 5188 7021 5216
rect 6788 5176 6794 5188
rect 7009 5185 7021 5188
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 11514 5216 11520 5228
rect 7156 5188 11520 5216
rect 7156 5176 7162 5188
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 2590 5148 2596 5160
rect 2551 5120 2596 5148
rect 2590 5108 2596 5120
rect 2648 5108 2654 5160
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5148 4399 5151
rect 4522 5148 4528 5160
rect 4387 5120 4528 5148
rect 4387 5117 4399 5120
rect 4341 5111 4399 5117
rect 4522 5108 4528 5120
rect 4580 5148 4586 5160
rect 5902 5148 5908 5160
rect 4580 5120 5908 5148
rect 4580 5108 4586 5120
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 8110 5148 8116 5160
rect 6052 5120 8116 5148
rect 6052 5108 6058 5120
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 4062 5040 4068 5092
rect 4120 5080 4126 5092
rect 6730 5080 6736 5092
rect 4120 5052 6736 5080
rect 4120 5040 4126 5052
rect 6730 5040 6736 5052
rect 6788 5040 6794 5092
rect 7193 5083 7251 5089
rect 7193 5049 7205 5083
rect 7239 5080 7251 5083
rect 7282 5080 7288 5092
rect 7239 5052 7288 5080
rect 7239 5049 7251 5052
rect 7193 5043 7251 5049
rect 7282 5040 7288 5052
rect 7340 5080 7346 5092
rect 11790 5080 11796 5092
rect 7340 5052 11796 5080
rect 7340 5040 7346 5052
rect 11790 5040 11796 5052
rect 11848 5040 11854 5092
rect 4617 5015 4675 5021
rect 4617 4981 4629 5015
rect 4663 5012 4675 5015
rect 4706 5012 4712 5024
rect 4663 4984 4712 5012
rect 4663 4981 4675 4984
rect 4617 4975 4675 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 4798 4972 4804 5024
rect 4856 5012 4862 5024
rect 5261 5015 5319 5021
rect 5261 5012 5273 5015
rect 4856 4984 5273 5012
rect 4856 4972 4862 4984
rect 5261 4981 5273 4984
rect 5307 4981 5319 5015
rect 5261 4975 5319 4981
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 6178 5012 6184 5024
rect 5408 4984 6184 5012
rect 5408 4972 5414 4984
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 8202 5012 8208 5024
rect 6420 4984 8208 5012
rect 6420 4972 6426 4984
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 1104 4922 16836 4944
rect 1104 4870 2924 4922
rect 2976 4870 2988 4922
rect 3040 4870 3052 4922
rect 3104 4870 3116 4922
rect 3168 4870 3180 4922
rect 3232 4870 6872 4922
rect 6924 4870 6936 4922
rect 6988 4870 7000 4922
rect 7052 4870 7064 4922
rect 7116 4870 7128 4922
rect 7180 4870 10820 4922
rect 10872 4870 10884 4922
rect 10936 4870 10948 4922
rect 11000 4870 11012 4922
rect 11064 4870 11076 4922
rect 11128 4870 14768 4922
rect 14820 4870 14832 4922
rect 14884 4870 14896 4922
rect 14948 4870 14960 4922
rect 15012 4870 15024 4922
rect 15076 4870 16836 4922
rect 1104 4848 16836 4870
rect 3050 4808 3056 4820
rect 3011 4780 3056 4808
rect 3050 4768 3056 4780
rect 3108 4768 3114 4820
rect 4062 4808 4068 4820
rect 3160 4780 4068 4808
rect 2685 4743 2743 4749
rect 2685 4709 2697 4743
rect 2731 4740 2743 4743
rect 3160 4740 3188 4780
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 4249 4811 4307 4817
rect 4249 4777 4261 4811
rect 4295 4808 4307 4811
rect 4522 4808 4528 4820
rect 4295 4780 4528 4808
rect 4295 4777 4307 4780
rect 4249 4771 4307 4777
rect 4522 4768 4528 4780
rect 4580 4808 4586 4820
rect 4580 4780 5764 4808
rect 4580 4768 4586 4780
rect 2731 4712 3188 4740
rect 3237 4743 3295 4749
rect 2731 4709 2743 4712
rect 2685 4703 2743 4709
rect 3237 4709 3249 4743
rect 3283 4740 3295 4743
rect 5534 4740 5540 4752
rect 3283 4712 5540 4740
rect 3283 4709 3295 4712
rect 3237 4703 3295 4709
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 5736 4740 5764 4780
rect 5810 4768 5816 4820
rect 5868 4808 5874 4820
rect 6089 4811 6147 4817
rect 6089 4808 6101 4811
rect 5868 4780 6101 4808
rect 5868 4768 5874 4780
rect 6089 4777 6101 4780
rect 6135 4777 6147 4811
rect 6089 4771 6147 4777
rect 6178 4768 6184 4820
rect 6236 4808 6242 4820
rect 6236 4780 6684 4808
rect 6236 4768 6242 4780
rect 6546 4740 6552 4752
rect 5736 4712 6552 4740
rect 6546 4700 6552 4712
rect 6604 4700 6610 4752
rect 6656 4740 6684 4780
rect 6730 4768 6736 4820
rect 6788 4808 6794 4820
rect 6825 4811 6883 4817
rect 6825 4808 6837 4811
rect 6788 4780 6837 4808
rect 6788 4768 6794 4780
rect 6825 4777 6837 4780
rect 6871 4777 6883 4811
rect 6825 4771 6883 4777
rect 9490 4740 9496 4752
rect 6656 4712 9496 4740
rect 9490 4700 9496 4712
rect 9548 4700 9554 4752
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 1670 4672 1676 4684
rect 1631 4644 1676 4672
rect 1670 4632 1676 4644
rect 1728 4632 1734 4684
rect 4430 4672 4436 4684
rect 3804 4644 4436 4672
rect 2682 4564 2688 4616
rect 2740 4604 2746 4616
rect 3804 4613 3832 4644
rect 4430 4632 4436 4644
rect 4488 4632 4494 4684
rect 4982 4672 4988 4684
rect 4540 4644 4988 4672
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 2740 4576 3801 4604
rect 2740 4564 2746 4576
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 4062 4604 4068 4616
rect 3975 4576 4068 4604
rect 3789 4567 3847 4573
rect 4062 4564 4068 4576
rect 4120 4604 4126 4616
rect 4540 4604 4568 4644
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 5445 4675 5503 4681
rect 5445 4641 5457 4675
rect 5491 4672 5503 4675
rect 7190 4672 7196 4684
rect 5491 4644 7196 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 4120 4576 4568 4604
rect 4120 4564 4126 4576
rect 4614 4564 4620 4616
rect 4672 4604 4678 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4672 4576 4721 4604
rect 4672 4564 4678 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 5353 4607 5411 4613
rect 5353 4606 5365 4607
rect 5276 4604 5365 4606
rect 4709 4567 4767 4573
rect 4816 4578 5365 4604
rect 4816 4576 5304 4578
rect 3881 4539 3939 4545
rect 3881 4536 3893 4539
rect 2746 4508 3893 4536
rect 2222 4428 2228 4480
rect 2280 4468 2286 4480
rect 2746 4468 2774 4508
rect 3881 4505 3893 4508
rect 3927 4505 3939 4539
rect 3881 4499 3939 4505
rect 4338 4496 4344 4548
rect 4396 4536 4402 4548
rect 4816 4536 4844 4576
rect 5353 4573 5365 4578
rect 5399 4573 5411 4607
rect 5994 4604 6000 4616
rect 5955 4576 6000 4604
rect 5353 4567 5411 4573
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 6178 4604 6184 4616
rect 6139 4576 6184 4604
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 6638 4604 6644 4616
rect 6599 4576 6644 4604
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 4396 4508 4844 4536
rect 4396 4496 4402 4508
rect 4982 4496 4988 4548
rect 5040 4536 5046 4548
rect 6196 4536 6224 4564
rect 12434 4536 12440 4548
rect 5040 4508 5488 4536
rect 6196 4508 12440 4536
rect 5040 4496 5046 4508
rect 2280 4440 2774 4468
rect 3053 4471 3111 4477
rect 2280 4428 2286 4440
rect 3053 4437 3065 4471
rect 3099 4468 3111 4471
rect 4154 4468 4160 4480
rect 3099 4440 4160 4468
rect 3099 4437 3111 4440
rect 3053 4431 3111 4437
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 4893 4471 4951 4477
rect 4893 4437 4905 4471
rect 4939 4468 4951 4471
rect 5350 4468 5356 4480
rect 4939 4440 5356 4468
rect 4939 4437 4951 4440
rect 4893 4431 4951 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 5460 4468 5488 4508
rect 12434 4496 12440 4508
rect 12492 4496 12498 4548
rect 9858 4468 9864 4480
rect 5460 4440 9864 4468
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 1104 4378 16836 4400
rect 1104 4326 4898 4378
rect 4950 4326 4962 4378
rect 5014 4326 5026 4378
rect 5078 4326 5090 4378
rect 5142 4326 5154 4378
rect 5206 4326 8846 4378
rect 8898 4326 8910 4378
rect 8962 4326 8974 4378
rect 9026 4326 9038 4378
rect 9090 4326 9102 4378
rect 9154 4326 12794 4378
rect 12846 4326 12858 4378
rect 12910 4326 12922 4378
rect 12974 4326 12986 4378
rect 13038 4326 13050 4378
rect 13102 4326 16836 4378
rect 1104 4304 16836 4326
rect 2685 4267 2743 4273
rect 2685 4233 2697 4267
rect 2731 4264 2743 4267
rect 2866 4264 2872 4276
rect 2731 4236 2872 4264
rect 2731 4233 2743 4236
rect 2685 4227 2743 4233
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 7742 4264 7748 4276
rect 3016 4236 7748 4264
rect 3016 4224 3022 4236
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 3602 4196 3608 4208
rect 3563 4168 3608 4196
rect 3602 4156 3608 4168
rect 3660 4156 3666 4208
rect 3789 4199 3847 4205
rect 3789 4165 3801 4199
rect 3835 4196 3847 4199
rect 4246 4196 4252 4208
rect 3835 4168 4252 4196
rect 3835 4165 3847 4168
rect 3789 4159 3847 4165
rect 4246 4156 4252 4168
rect 4304 4156 4310 4208
rect 4522 4196 4528 4208
rect 4448 4168 4528 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 1762 4128 1768 4140
rect 1719 4100 1768 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 1762 4088 1768 4100
rect 1820 4088 1826 4140
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 3053 4131 3111 4137
rect 2924 4100 2969 4128
rect 2924 4088 2930 4100
rect 3053 4097 3065 4131
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 4448 4128 4476 4168
rect 4522 4156 4528 4168
rect 4580 4156 4586 4208
rect 5994 4196 6000 4208
rect 5092 4168 6000 4196
rect 5092 4140 5120 4168
rect 5994 4156 6000 4168
rect 6052 4156 6058 4208
rect 4614 4128 4620 4140
rect 3191 4100 4476 4128
rect 4575 4100 4620 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 1394 4060 1400 4072
rect 1355 4032 1400 4060
rect 1394 4020 1400 4032
rect 1452 4020 1458 4072
rect 2498 4020 2504 4072
rect 2556 4060 2562 4072
rect 2958 4060 2964 4072
rect 2556 4032 2964 4060
rect 2556 4020 2562 4032
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3068 3924 3096 4091
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 5074 4128 5080 4140
rect 4987 4100 5080 4128
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4128 5319 4131
rect 6178 4128 6184 4140
rect 5307 4100 6184 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 3970 4060 3976 4072
rect 3931 4032 3976 4060
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 5276 4060 5304 4091
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 5092 4032 5304 4060
rect 3878 3952 3884 4004
rect 3936 3992 3942 4004
rect 5092 3992 5120 4032
rect 3936 3964 5120 3992
rect 5169 3995 5227 4001
rect 3936 3952 3942 3964
rect 5169 3961 5181 3995
rect 5215 3992 5227 3995
rect 5258 3992 5264 4004
rect 5215 3964 5264 3992
rect 5215 3961 5227 3964
rect 5169 3955 5227 3961
rect 5258 3952 5264 3964
rect 5316 3952 5322 4004
rect 4338 3924 4344 3936
rect 3068 3896 4344 3924
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 7374 3924 7380 3936
rect 4571 3896 7380 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 1104 3834 16836 3856
rect 1104 3782 2924 3834
rect 2976 3782 2988 3834
rect 3040 3782 3052 3834
rect 3104 3782 3116 3834
rect 3168 3782 3180 3834
rect 3232 3782 6872 3834
rect 6924 3782 6936 3834
rect 6988 3782 7000 3834
rect 7052 3782 7064 3834
rect 7116 3782 7128 3834
rect 7180 3782 10820 3834
rect 10872 3782 10884 3834
rect 10936 3782 10948 3834
rect 11000 3782 11012 3834
rect 11064 3782 11076 3834
rect 11128 3782 14768 3834
rect 14820 3782 14832 3834
rect 14884 3782 14896 3834
rect 14948 3782 14960 3834
rect 15012 3782 15024 3834
rect 15076 3782 16836 3834
rect 1104 3760 16836 3782
rect 2314 3680 2320 3732
rect 2372 3720 2378 3732
rect 3881 3723 3939 3729
rect 3881 3720 3893 3723
rect 2372 3692 3893 3720
rect 2372 3680 2378 3692
rect 3881 3689 3893 3692
rect 3927 3689 3939 3723
rect 3881 3683 3939 3689
rect 4338 3680 4344 3732
rect 4396 3720 4402 3732
rect 11238 3720 11244 3732
rect 4396 3692 11244 3720
rect 4396 3680 4402 3692
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 2682 3652 2688 3664
rect 2148 3624 2688 3652
rect 2038 3584 2044 3596
rect 1504 3556 2044 3584
rect 1504 3525 1532 3556
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3485 1547 3519
rect 1670 3516 1676 3528
rect 1631 3488 1676 3516
rect 1489 3479 1547 3485
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 2148 3525 2176 3624
rect 2682 3612 2688 3624
rect 2740 3612 2746 3664
rect 3053 3655 3111 3661
rect 3053 3621 3065 3655
rect 3099 3621 3111 3655
rect 3053 3615 3111 3621
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3584 2375 3587
rect 2363 3556 2452 3584
rect 2363 3553 2375 3556
rect 2317 3547 2375 3553
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2222 3476 2228 3528
rect 2280 3516 2286 3528
rect 2280 3488 2325 3516
rect 2280 3476 2286 3488
rect 1581 3451 1639 3457
rect 1581 3417 1593 3451
rect 1627 3448 1639 3451
rect 2240 3448 2268 3476
rect 1627 3420 2268 3448
rect 2424 3448 2452 3556
rect 3068 3528 3096 3615
rect 3694 3612 3700 3664
rect 3752 3652 3758 3664
rect 4433 3655 4491 3661
rect 4433 3652 4445 3655
rect 3752 3624 4445 3652
rect 3752 3612 3758 3624
rect 4433 3621 4445 3624
rect 4479 3621 4491 3655
rect 4433 3615 4491 3621
rect 5074 3584 5080 3596
rect 3988 3556 5080 3584
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 2958 3516 2964 3528
rect 2547 3488 2887 3516
rect 2919 3488 2964 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 2859 3448 2887 3488
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3050 3476 3056 3528
rect 3108 3476 3114 3528
rect 3142 3476 3148 3528
rect 3200 3516 3206 3528
rect 3789 3519 3847 3525
rect 3200 3488 3245 3516
rect 3200 3476 3206 3488
rect 3789 3485 3801 3519
rect 3835 3516 3847 3519
rect 3878 3516 3884 3528
rect 3835 3488 3884 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 3988 3525 4016 3556
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 8294 3516 8300 3528
rect 4663 3488 8300 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 11330 3448 11336 3460
rect 2424 3420 2544 3448
rect 2859 3420 11336 3448
rect 1627 3417 1639 3420
rect 1581 3411 1639 3417
rect 2130 3340 2136 3392
rect 2188 3380 2194 3392
rect 2409 3383 2467 3389
rect 2409 3380 2421 3383
rect 2188 3352 2421 3380
rect 2188 3340 2194 3352
rect 2409 3349 2421 3352
rect 2455 3349 2467 3383
rect 2516 3380 2544 3420
rect 11330 3408 11336 3420
rect 11388 3408 11394 3460
rect 4062 3380 4068 3392
rect 2516 3352 4068 3380
rect 2409 3343 2467 3349
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 1104 3290 16836 3312
rect 1104 3238 4898 3290
rect 4950 3238 4962 3290
rect 5014 3238 5026 3290
rect 5078 3238 5090 3290
rect 5142 3238 5154 3290
rect 5206 3238 8846 3290
rect 8898 3238 8910 3290
rect 8962 3238 8974 3290
rect 9026 3238 9038 3290
rect 9090 3238 9102 3290
rect 9154 3238 12794 3290
rect 12846 3238 12858 3290
rect 12910 3238 12922 3290
rect 12974 3238 12986 3290
rect 13038 3238 13050 3290
rect 13102 3238 16836 3290
rect 1104 3216 16836 3238
rect 2406 3176 2412 3188
rect 2367 3148 2412 3176
rect 2406 3136 2412 3148
rect 2464 3136 2470 3188
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3326 3176 3332 3188
rect 3099 3148 3332 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 1854 3068 1860 3120
rect 1912 3108 1918 3120
rect 3142 3108 3148 3120
rect 1912 3080 3148 3108
rect 1912 3068 1918 3080
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 1489 3043 1547 3049
rect 1489 3009 1501 3043
rect 1535 3040 1547 3043
rect 1578 3040 1584 3052
rect 1535 3012 1584 3040
rect 1535 3009 1547 3012
rect 1489 3003 1547 3009
rect 1578 3000 1584 3012
rect 1636 3000 1642 3052
rect 2222 3040 2228 3052
rect 2183 3012 2228 3040
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 2556 3012 2881 3040
rect 2556 3000 2562 3012
rect 2869 3009 2881 3012
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 7926 3040 7932 3052
rect 3743 3012 7932 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 3068 2972 3096 3003
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 8386 2972 8392 2984
rect 3068 2944 8392 2972
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 3142 2864 3148 2916
rect 3200 2904 3206 2916
rect 3513 2907 3571 2913
rect 3513 2904 3525 2907
rect 3200 2876 3525 2904
rect 3200 2864 3206 2876
rect 3513 2873 3525 2876
rect 3559 2873 3571 2907
rect 3513 2867 3571 2873
rect 1673 2839 1731 2845
rect 1673 2805 1685 2839
rect 1719 2836 1731 2839
rect 9766 2836 9772 2848
rect 1719 2808 9772 2836
rect 1719 2805 1731 2808
rect 1673 2799 1731 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 1104 2746 16836 2768
rect 1104 2694 2924 2746
rect 2976 2694 2988 2746
rect 3040 2694 3052 2746
rect 3104 2694 3116 2746
rect 3168 2694 3180 2746
rect 3232 2694 6872 2746
rect 6924 2694 6936 2746
rect 6988 2694 7000 2746
rect 7052 2694 7064 2746
rect 7116 2694 7128 2746
rect 7180 2694 10820 2746
rect 10872 2694 10884 2746
rect 10936 2694 10948 2746
rect 11000 2694 11012 2746
rect 11064 2694 11076 2746
rect 11128 2694 14768 2746
rect 14820 2694 14832 2746
rect 14884 2694 14896 2746
rect 14948 2694 14960 2746
rect 15012 2694 15024 2746
rect 15076 2694 16836 2746
rect 1104 2672 16836 2694
rect 1946 2592 1952 2644
rect 2004 2632 2010 2644
rect 2869 2635 2927 2641
rect 2869 2632 2881 2635
rect 2004 2604 2881 2632
rect 2004 2592 2010 2604
rect 2869 2601 2881 2604
rect 2915 2601 2927 2635
rect 2869 2595 2927 2601
rect 2682 2524 2688 2576
rect 2740 2524 2746 2576
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 2038 2496 2044 2508
rect 1719 2468 2044 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 2038 2456 2044 2468
rect 2096 2496 2102 2508
rect 2700 2496 2728 2524
rect 2096 2468 2728 2496
rect 2096 2456 2102 2468
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 2682 2428 2688 2440
rect 2643 2400 2688 2428
rect 2682 2388 2688 2400
rect 2740 2428 2746 2440
rect 5718 2428 5724 2440
rect 2740 2400 5724 2428
rect 2740 2388 2746 2400
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 1104 2202 16836 2224
rect 1104 2150 4898 2202
rect 4950 2150 4962 2202
rect 5014 2150 5026 2202
rect 5078 2150 5090 2202
rect 5142 2150 5154 2202
rect 5206 2150 8846 2202
rect 8898 2150 8910 2202
rect 8962 2150 8974 2202
rect 9026 2150 9038 2202
rect 9090 2150 9102 2202
rect 9154 2150 12794 2202
rect 12846 2150 12858 2202
rect 12910 2150 12922 2202
rect 12974 2150 12986 2202
rect 13038 2150 13050 2202
rect 13102 2150 16836 2202
rect 1104 2128 16836 2150
rect 1581 2091 1639 2097
rect 1581 2057 1593 2091
rect 1627 2088 1639 2091
rect 3602 2088 3608 2100
rect 1627 2060 3608 2088
rect 1627 2057 1639 2060
rect 1581 2051 1639 2057
rect 3602 2048 3608 2060
rect 3660 2048 3666 2100
rect 3418 2020 3424 2032
rect 1412 1992 3424 2020
rect 1412 1961 1440 1992
rect 3418 1980 3424 1992
rect 3476 1980 3482 2032
rect 1397 1955 1455 1961
rect 1397 1921 1409 1955
rect 1443 1921 1455 1955
rect 2038 1952 2044 1964
rect 1999 1924 2044 1952
rect 1397 1915 1455 1921
rect 2038 1912 2044 1924
rect 2096 1912 2102 1964
rect 2225 1955 2283 1961
rect 2225 1921 2237 1955
rect 2271 1952 2283 1955
rect 2682 1952 2688 1964
rect 2271 1924 2688 1952
rect 2271 1921 2283 1924
rect 2225 1915 2283 1921
rect 2682 1912 2688 1924
rect 2740 1912 2746 1964
rect 2133 1887 2191 1893
rect 2133 1853 2145 1887
rect 2179 1884 2191 1887
rect 2774 1884 2780 1896
rect 2179 1856 2780 1884
rect 2179 1853 2191 1856
rect 2133 1847 2191 1853
rect 2774 1844 2780 1856
rect 2832 1844 2838 1896
rect 1104 1658 16836 1680
rect 1104 1606 2924 1658
rect 2976 1606 2988 1658
rect 3040 1606 3052 1658
rect 3104 1606 3116 1658
rect 3168 1606 3180 1658
rect 3232 1606 6872 1658
rect 6924 1606 6936 1658
rect 6988 1606 7000 1658
rect 7052 1606 7064 1658
rect 7116 1606 7128 1658
rect 7180 1606 10820 1658
rect 10872 1606 10884 1658
rect 10936 1606 10948 1658
rect 11000 1606 11012 1658
rect 11064 1606 11076 1658
rect 11128 1606 14768 1658
rect 14820 1606 14832 1658
rect 14884 1606 14896 1658
rect 14948 1606 14960 1658
rect 15012 1606 15024 1658
rect 15076 1606 16836 1658
rect 1104 1584 16836 1606
rect 1394 1340 1400 1352
rect 1355 1312 1400 1340
rect 1394 1300 1400 1312
rect 1452 1300 1458 1352
rect 1486 1164 1492 1216
rect 1544 1204 1550 1216
rect 1581 1207 1639 1213
rect 1581 1204 1593 1207
rect 1544 1176 1593 1204
rect 1544 1164 1550 1176
rect 1581 1173 1593 1176
rect 1627 1173 1639 1207
rect 1581 1167 1639 1173
rect 1104 1114 16836 1136
rect 1104 1062 4898 1114
rect 4950 1062 4962 1114
rect 5014 1062 5026 1114
rect 5078 1062 5090 1114
rect 5142 1062 5154 1114
rect 5206 1062 8846 1114
rect 8898 1062 8910 1114
rect 8962 1062 8974 1114
rect 9026 1062 9038 1114
rect 9090 1062 9102 1114
rect 9154 1062 12794 1114
rect 12846 1062 12858 1114
rect 12910 1062 12922 1114
rect 12974 1062 12986 1114
rect 13038 1062 13050 1114
rect 13102 1062 16836 1114
rect 1104 1040 16836 1062
<< via1 >>
rect 4898 22822 4950 22874
rect 4962 22822 5014 22874
rect 5026 22822 5078 22874
rect 5090 22822 5142 22874
rect 5154 22822 5206 22874
rect 8846 22822 8898 22874
rect 8910 22822 8962 22874
rect 8974 22822 9026 22874
rect 9038 22822 9090 22874
rect 9102 22822 9154 22874
rect 12794 22822 12846 22874
rect 12858 22822 12910 22874
rect 12922 22822 12974 22874
rect 12986 22822 13038 22874
rect 13050 22822 13102 22874
rect 2924 22278 2976 22330
rect 2988 22278 3040 22330
rect 3052 22278 3104 22330
rect 3116 22278 3168 22330
rect 3180 22278 3232 22330
rect 6872 22278 6924 22330
rect 6936 22278 6988 22330
rect 7000 22278 7052 22330
rect 7064 22278 7116 22330
rect 7128 22278 7180 22330
rect 10820 22278 10872 22330
rect 10884 22278 10936 22330
rect 10948 22278 11000 22330
rect 11012 22278 11064 22330
rect 11076 22278 11128 22330
rect 14768 22278 14820 22330
rect 14832 22278 14884 22330
rect 14896 22278 14948 22330
rect 14960 22278 15012 22330
rect 15024 22278 15076 22330
rect 4898 21734 4950 21786
rect 4962 21734 5014 21786
rect 5026 21734 5078 21786
rect 5090 21734 5142 21786
rect 5154 21734 5206 21786
rect 8846 21734 8898 21786
rect 8910 21734 8962 21786
rect 8974 21734 9026 21786
rect 9038 21734 9090 21786
rect 9102 21734 9154 21786
rect 12794 21734 12846 21786
rect 12858 21734 12910 21786
rect 12922 21734 12974 21786
rect 12986 21734 13038 21786
rect 13050 21734 13102 21786
rect 2924 21190 2976 21242
rect 2988 21190 3040 21242
rect 3052 21190 3104 21242
rect 3116 21190 3168 21242
rect 3180 21190 3232 21242
rect 6872 21190 6924 21242
rect 6936 21190 6988 21242
rect 7000 21190 7052 21242
rect 7064 21190 7116 21242
rect 7128 21190 7180 21242
rect 10820 21190 10872 21242
rect 10884 21190 10936 21242
rect 10948 21190 11000 21242
rect 11012 21190 11064 21242
rect 11076 21190 11128 21242
rect 14768 21190 14820 21242
rect 14832 21190 14884 21242
rect 14896 21190 14948 21242
rect 14960 21190 15012 21242
rect 15024 21190 15076 21242
rect 4898 20646 4950 20698
rect 4962 20646 5014 20698
rect 5026 20646 5078 20698
rect 5090 20646 5142 20698
rect 5154 20646 5206 20698
rect 8846 20646 8898 20698
rect 8910 20646 8962 20698
rect 8974 20646 9026 20698
rect 9038 20646 9090 20698
rect 9102 20646 9154 20698
rect 12794 20646 12846 20698
rect 12858 20646 12910 20698
rect 12922 20646 12974 20698
rect 12986 20646 13038 20698
rect 13050 20646 13102 20698
rect 2780 20544 2832 20596
rect 1676 20451 1728 20460
rect 1676 20417 1685 20451
rect 1685 20417 1719 20451
rect 1719 20417 1728 20451
rect 1676 20408 1728 20417
rect 2924 20102 2976 20154
rect 2988 20102 3040 20154
rect 3052 20102 3104 20154
rect 3116 20102 3168 20154
rect 3180 20102 3232 20154
rect 6872 20102 6924 20154
rect 6936 20102 6988 20154
rect 7000 20102 7052 20154
rect 7064 20102 7116 20154
rect 7128 20102 7180 20154
rect 10820 20102 10872 20154
rect 10884 20102 10936 20154
rect 10948 20102 11000 20154
rect 11012 20102 11064 20154
rect 11076 20102 11128 20154
rect 14768 20102 14820 20154
rect 14832 20102 14884 20154
rect 14896 20102 14948 20154
rect 14960 20102 15012 20154
rect 15024 20102 15076 20154
rect 4898 19558 4950 19610
rect 4962 19558 5014 19610
rect 5026 19558 5078 19610
rect 5090 19558 5142 19610
rect 5154 19558 5206 19610
rect 8846 19558 8898 19610
rect 8910 19558 8962 19610
rect 8974 19558 9026 19610
rect 9038 19558 9090 19610
rect 9102 19558 9154 19610
rect 12794 19558 12846 19610
rect 12858 19558 12910 19610
rect 12922 19558 12974 19610
rect 12986 19558 13038 19610
rect 13050 19558 13102 19610
rect 2924 19014 2976 19066
rect 2988 19014 3040 19066
rect 3052 19014 3104 19066
rect 3116 19014 3168 19066
rect 3180 19014 3232 19066
rect 6872 19014 6924 19066
rect 6936 19014 6988 19066
rect 7000 19014 7052 19066
rect 7064 19014 7116 19066
rect 7128 19014 7180 19066
rect 10820 19014 10872 19066
rect 10884 19014 10936 19066
rect 10948 19014 11000 19066
rect 11012 19014 11064 19066
rect 11076 19014 11128 19066
rect 14768 19014 14820 19066
rect 14832 19014 14884 19066
rect 14896 19014 14948 19066
rect 14960 19014 15012 19066
rect 15024 19014 15076 19066
rect 1492 18955 1544 18964
rect 1492 18921 1501 18955
rect 1501 18921 1535 18955
rect 1535 18921 1544 18955
rect 1492 18912 1544 18921
rect 1676 18912 1728 18964
rect 2320 18751 2372 18760
rect 2320 18717 2329 18751
rect 2329 18717 2363 18751
rect 2363 18717 2372 18751
rect 2320 18708 2372 18717
rect 4804 18640 4856 18692
rect 4898 18470 4950 18522
rect 4962 18470 5014 18522
rect 5026 18470 5078 18522
rect 5090 18470 5142 18522
rect 5154 18470 5206 18522
rect 8846 18470 8898 18522
rect 8910 18470 8962 18522
rect 8974 18470 9026 18522
rect 9038 18470 9090 18522
rect 9102 18470 9154 18522
rect 12794 18470 12846 18522
rect 12858 18470 12910 18522
rect 12922 18470 12974 18522
rect 12986 18470 13038 18522
rect 13050 18470 13102 18522
rect 2412 18232 2464 18284
rect 3700 18164 3752 18216
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 2136 18071 2188 18080
rect 2136 18037 2145 18071
rect 2145 18037 2179 18071
rect 2179 18037 2188 18071
rect 2136 18028 2188 18037
rect 2924 17926 2976 17978
rect 2988 17926 3040 17978
rect 3052 17926 3104 17978
rect 3116 17926 3168 17978
rect 3180 17926 3232 17978
rect 6872 17926 6924 17978
rect 6936 17926 6988 17978
rect 7000 17926 7052 17978
rect 7064 17926 7116 17978
rect 7128 17926 7180 17978
rect 10820 17926 10872 17978
rect 10884 17926 10936 17978
rect 10948 17926 11000 17978
rect 11012 17926 11064 17978
rect 11076 17926 11128 17978
rect 14768 17926 14820 17978
rect 14832 17926 14884 17978
rect 14896 17926 14948 17978
rect 14960 17926 15012 17978
rect 15024 17926 15076 17978
rect 2780 17824 2832 17876
rect 3332 17824 3384 17876
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 4528 17620 4580 17672
rect 3332 17552 3384 17604
rect 4898 17382 4950 17434
rect 4962 17382 5014 17434
rect 5026 17382 5078 17434
rect 5090 17382 5142 17434
rect 5154 17382 5206 17434
rect 8846 17382 8898 17434
rect 8910 17382 8962 17434
rect 8974 17382 9026 17434
rect 9038 17382 9090 17434
rect 9102 17382 9154 17434
rect 12794 17382 12846 17434
rect 12858 17382 12910 17434
rect 12922 17382 12974 17434
rect 12986 17382 13038 17434
rect 13050 17382 13102 17434
rect 2320 17280 2372 17332
rect 3700 17323 3752 17332
rect 3700 17289 3709 17323
rect 3709 17289 3743 17323
rect 3743 17289 3752 17323
rect 3700 17280 3752 17289
rect 11336 17212 11388 17264
rect 1492 17076 1544 17128
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 2320 17076 2372 17128
rect 6276 17008 6328 17060
rect 3516 16940 3568 16992
rect 2924 16838 2976 16890
rect 2988 16838 3040 16890
rect 3052 16838 3104 16890
rect 3116 16838 3168 16890
rect 3180 16838 3232 16890
rect 6872 16838 6924 16890
rect 6936 16838 6988 16890
rect 7000 16838 7052 16890
rect 7064 16838 7116 16890
rect 7128 16838 7180 16890
rect 10820 16838 10872 16890
rect 10884 16838 10936 16890
rect 10948 16838 11000 16890
rect 11012 16838 11064 16890
rect 11076 16838 11128 16890
rect 14768 16838 14820 16890
rect 14832 16838 14884 16890
rect 14896 16838 14948 16890
rect 14960 16838 15012 16890
rect 15024 16838 15076 16890
rect 1952 16668 2004 16720
rect 4344 16668 4396 16720
rect 9220 16600 9272 16652
rect 4712 16575 4764 16584
rect 2504 16464 2556 16516
rect 3056 16507 3108 16516
rect 3056 16473 3065 16507
rect 3065 16473 3099 16507
rect 3099 16473 3108 16507
rect 3056 16464 3108 16473
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 4712 16532 4764 16541
rect 1952 16439 2004 16448
rect 1952 16405 1961 16439
rect 1961 16405 1995 16439
rect 1995 16405 2004 16439
rect 1952 16396 2004 16405
rect 2044 16439 2096 16448
rect 2044 16405 2053 16439
rect 2053 16405 2087 16439
rect 2087 16405 2096 16439
rect 2412 16439 2464 16448
rect 2044 16396 2096 16405
rect 2412 16405 2421 16439
rect 2421 16405 2455 16439
rect 2455 16405 2464 16439
rect 2412 16396 2464 16405
rect 2780 16396 2832 16448
rect 6736 16464 6788 16516
rect 3976 16396 4028 16448
rect 4898 16294 4950 16346
rect 4962 16294 5014 16346
rect 5026 16294 5078 16346
rect 5090 16294 5142 16346
rect 5154 16294 5206 16346
rect 8846 16294 8898 16346
rect 8910 16294 8962 16346
rect 8974 16294 9026 16346
rect 9038 16294 9090 16346
rect 9102 16294 9154 16346
rect 12794 16294 12846 16346
rect 12858 16294 12910 16346
rect 12922 16294 12974 16346
rect 12986 16294 13038 16346
rect 13050 16294 13102 16346
rect 4528 16235 4580 16244
rect 4528 16201 4537 16235
rect 4537 16201 4571 16235
rect 4571 16201 4580 16235
rect 4528 16192 4580 16201
rect 1676 16056 1728 16108
rect 5448 16056 5500 16108
rect 5816 16099 5868 16108
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 3424 15988 3476 16040
rect 3608 15988 3660 16040
rect 3884 15988 3936 16040
rect 4344 15988 4396 16040
rect 7932 15920 7984 15972
rect 2136 15852 2188 15904
rect 3056 15852 3108 15904
rect 5264 15852 5316 15904
rect 6092 15852 6144 15904
rect 2924 15750 2976 15802
rect 2988 15750 3040 15802
rect 3052 15750 3104 15802
rect 3116 15750 3168 15802
rect 3180 15750 3232 15802
rect 6872 15750 6924 15802
rect 6936 15750 6988 15802
rect 7000 15750 7052 15802
rect 7064 15750 7116 15802
rect 7128 15750 7180 15802
rect 10820 15750 10872 15802
rect 10884 15750 10936 15802
rect 10948 15750 11000 15802
rect 11012 15750 11064 15802
rect 11076 15750 11128 15802
rect 14768 15750 14820 15802
rect 14832 15750 14884 15802
rect 14896 15750 14948 15802
rect 14960 15750 15012 15802
rect 15024 15750 15076 15802
rect 4804 15648 4856 15700
rect 5264 15648 5316 15700
rect 9588 15648 9640 15700
rect 6460 15580 6512 15632
rect 4160 15512 4212 15564
rect 5724 15512 5776 15564
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 4344 15487 4396 15496
rect 4344 15453 4353 15487
rect 4353 15453 4387 15487
rect 4387 15453 4396 15487
rect 4344 15444 4396 15453
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 4068 15376 4120 15428
rect 6184 15444 6236 15496
rect 7380 15444 7432 15496
rect 3608 15308 3660 15360
rect 7196 15376 7248 15428
rect 5816 15308 5868 15360
rect 4898 15206 4950 15258
rect 4962 15206 5014 15258
rect 5026 15206 5078 15258
rect 5090 15206 5142 15258
rect 5154 15206 5206 15258
rect 8846 15206 8898 15258
rect 8910 15206 8962 15258
rect 8974 15206 9026 15258
rect 9038 15206 9090 15258
rect 9102 15206 9154 15258
rect 12794 15206 12846 15258
rect 12858 15206 12910 15258
rect 12922 15206 12974 15258
rect 12986 15206 13038 15258
rect 13050 15206 13102 15258
rect 8484 15104 8536 15156
rect 4068 15036 4120 15088
rect 8576 15036 8628 15088
rect 4252 14968 4304 15020
rect 5724 15011 5776 15020
rect 5724 14977 5733 15011
rect 5733 14977 5767 15011
rect 5767 14977 5776 15011
rect 5724 14968 5776 14977
rect 6000 14968 6052 15020
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 3424 14900 3476 14952
rect 5356 14900 5408 14952
rect 7012 14968 7064 15020
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 8760 14900 8812 14952
rect 6368 14875 6420 14884
rect 6368 14841 6377 14875
rect 6377 14841 6411 14875
rect 6411 14841 6420 14875
rect 6368 14832 6420 14841
rect 7012 14832 7064 14884
rect 8392 14832 8444 14884
rect 4528 14764 4580 14816
rect 4620 14764 4672 14816
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 8300 14764 8352 14816
rect 2924 14662 2976 14714
rect 2988 14662 3040 14714
rect 3052 14662 3104 14714
rect 3116 14662 3168 14714
rect 3180 14662 3232 14714
rect 6872 14662 6924 14714
rect 6936 14662 6988 14714
rect 7000 14662 7052 14714
rect 7064 14662 7116 14714
rect 7128 14662 7180 14714
rect 10820 14662 10872 14714
rect 10884 14662 10936 14714
rect 10948 14662 11000 14714
rect 11012 14662 11064 14714
rect 11076 14662 11128 14714
rect 14768 14662 14820 14714
rect 14832 14662 14884 14714
rect 14896 14662 14948 14714
rect 14960 14662 15012 14714
rect 15024 14662 15076 14714
rect 4160 14560 4212 14612
rect 4528 14560 4580 14612
rect 5448 14492 5500 14544
rect 6184 14560 6236 14612
rect 6552 14492 6604 14544
rect 6920 14424 6972 14476
rect 2228 14356 2280 14408
rect 7196 14424 7248 14476
rect 1676 14331 1728 14340
rect 1676 14297 1710 14331
rect 1710 14297 1728 14331
rect 1676 14288 1728 14297
rect 1768 14288 1820 14340
rect 2044 14288 2096 14340
rect 4436 14288 4488 14340
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 9312 14424 9364 14476
rect 3792 14263 3844 14272
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 7196 14288 7248 14340
rect 5816 14220 5868 14272
rect 6000 14263 6052 14272
rect 6000 14229 6009 14263
rect 6009 14229 6043 14263
rect 6043 14229 6052 14263
rect 6000 14220 6052 14229
rect 6368 14220 6420 14272
rect 7472 14220 7524 14272
rect 4898 14118 4950 14170
rect 4962 14118 5014 14170
rect 5026 14118 5078 14170
rect 5090 14118 5142 14170
rect 5154 14118 5206 14170
rect 8846 14118 8898 14170
rect 8910 14118 8962 14170
rect 8974 14118 9026 14170
rect 9038 14118 9090 14170
rect 9102 14118 9154 14170
rect 12794 14118 12846 14170
rect 12858 14118 12910 14170
rect 12922 14118 12974 14170
rect 12986 14118 13038 14170
rect 13050 14118 13102 14170
rect 6828 14016 6880 14068
rect 2044 13923 2096 13932
rect 2044 13889 2078 13923
rect 2078 13889 2096 13923
rect 2044 13880 2096 13889
rect 3976 13948 4028 14000
rect 4068 13948 4120 14000
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 5448 13812 5500 13864
rect 1676 13676 1728 13728
rect 5448 13676 5500 13728
rect 5908 13880 5960 13932
rect 7748 13923 7800 13932
rect 7748 13889 7757 13923
rect 7757 13889 7791 13923
rect 7791 13889 7800 13923
rect 7748 13880 7800 13889
rect 8208 13880 8260 13932
rect 8668 13923 8720 13932
rect 8668 13889 8677 13923
rect 8677 13889 8711 13923
rect 8711 13889 8720 13923
rect 8668 13880 8720 13889
rect 11612 13880 11664 13932
rect 5724 13812 5776 13864
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 8024 13855 8076 13864
rect 6920 13812 6972 13821
rect 5908 13744 5960 13796
rect 6276 13744 6328 13796
rect 6736 13744 6788 13796
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 9956 13812 10008 13864
rect 7196 13676 7248 13728
rect 2924 13574 2976 13626
rect 2988 13574 3040 13626
rect 3052 13574 3104 13626
rect 3116 13574 3168 13626
rect 3180 13574 3232 13626
rect 6872 13574 6924 13626
rect 6936 13574 6988 13626
rect 7000 13574 7052 13626
rect 7064 13574 7116 13626
rect 7128 13574 7180 13626
rect 10820 13574 10872 13626
rect 10884 13574 10936 13626
rect 10948 13574 11000 13626
rect 11012 13574 11064 13626
rect 11076 13574 11128 13626
rect 14768 13574 14820 13626
rect 14832 13574 14884 13626
rect 14896 13574 14948 13626
rect 14960 13574 15012 13626
rect 15024 13574 15076 13626
rect 6000 13472 6052 13524
rect 7288 13472 7340 13524
rect 9588 13472 9640 13524
rect 11060 13472 11112 13524
rect 7748 13404 7800 13456
rect 5448 13336 5500 13388
rect 3884 13268 3936 13320
rect 1768 13200 1820 13252
rect 2044 13200 2096 13252
rect 4252 13200 4304 13252
rect 3332 13132 3384 13184
rect 6460 13268 6512 13320
rect 7196 13268 7248 13320
rect 7564 13268 7616 13320
rect 6092 13200 6144 13252
rect 6552 13200 6604 13252
rect 6920 13200 6972 13252
rect 7288 13200 7340 13252
rect 8760 13336 8812 13388
rect 10692 13336 10744 13388
rect 8392 13268 8444 13320
rect 9864 13311 9916 13320
rect 9864 13277 9873 13311
rect 9873 13277 9907 13311
rect 9907 13277 9916 13311
rect 9864 13268 9916 13277
rect 8024 13132 8076 13184
rect 10508 13200 10560 13252
rect 11244 13132 11296 13184
rect 4898 13030 4950 13082
rect 4962 13030 5014 13082
rect 5026 13030 5078 13082
rect 5090 13030 5142 13082
rect 5154 13030 5206 13082
rect 8846 13030 8898 13082
rect 8910 13030 8962 13082
rect 8974 13030 9026 13082
rect 9038 13030 9090 13082
rect 9102 13030 9154 13082
rect 12794 13030 12846 13082
rect 12858 13030 12910 13082
rect 12922 13030 12974 13082
rect 12986 13030 13038 13082
rect 13050 13030 13102 13082
rect 1400 12971 1452 12980
rect 1400 12937 1409 12971
rect 1409 12937 1443 12971
rect 1443 12937 1452 12971
rect 1400 12928 1452 12937
rect 2228 12928 2280 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 6552 12928 6604 12980
rect 8300 12928 8352 12980
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 2688 12835 2740 12844
rect 2688 12801 2697 12835
rect 2697 12801 2731 12835
rect 2731 12801 2740 12835
rect 2964 12835 3016 12844
rect 2688 12792 2740 12801
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 3792 12792 3844 12844
rect 8024 12860 8076 12912
rect 9036 12860 9088 12912
rect 11980 12928 12032 12980
rect 4436 12792 4488 12844
rect 7656 12792 7708 12844
rect 8852 12792 8904 12844
rect 2320 12724 2372 12776
rect 3424 12656 3476 12708
rect 4160 12724 4212 12776
rect 8024 12724 8076 12776
rect 9680 12724 9732 12776
rect 8944 12656 8996 12708
rect 10048 12792 10100 12844
rect 11060 12792 11112 12844
rect 11428 12792 11480 12844
rect 7748 12588 7800 12640
rect 8392 12631 8444 12640
rect 8392 12597 8401 12631
rect 8401 12597 8435 12631
rect 8435 12597 8444 12631
rect 8392 12588 8444 12597
rect 8484 12588 8536 12640
rect 9220 12588 9272 12640
rect 9496 12588 9548 12640
rect 12164 12656 12216 12708
rect 10140 12588 10192 12640
rect 10232 12588 10284 12640
rect 11244 12588 11296 12640
rect 12072 12588 12124 12640
rect 2924 12486 2976 12538
rect 2988 12486 3040 12538
rect 3052 12486 3104 12538
rect 3116 12486 3168 12538
rect 3180 12486 3232 12538
rect 6872 12486 6924 12538
rect 6936 12486 6988 12538
rect 7000 12486 7052 12538
rect 7064 12486 7116 12538
rect 7128 12486 7180 12538
rect 10820 12486 10872 12538
rect 10884 12486 10936 12538
rect 10948 12486 11000 12538
rect 11012 12486 11064 12538
rect 11076 12486 11128 12538
rect 14768 12486 14820 12538
rect 14832 12486 14884 12538
rect 14896 12486 14948 12538
rect 14960 12486 15012 12538
rect 15024 12486 15076 12538
rect 2780 12384 2832 12436
rect 3976 12384 4028 12436
rect 7656 12384 7708 12436
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 8300 12427 8352 12436
rect 8300 12393 8309 12427
rect 8309 12393 8343 12427
rect 8343 12393 8352 12427
rect 8300 12384 8352 12393
rect 10416 12384 10468 12436
rect 10784 12427 10836 12436
rect 3056 12316 3108 12368
rect 3424 12316 3476 12368
rect 2136 12248 2188 12300
rect 2504 12248 2556 12300
rect 3332 12248 3384 12300
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 3792 12180 3844 12232
rect 4620 12291 4672 12300
rect 4620 12257 4638 12291
rect 4638 12257 4672 12291
rect 4620 12248 4672 12257
rect 4988 12291 5040 12300
rect 4988 12257 4997 12291
rect 4997 12257 5031 12291
rect 5031 12257 5040 12291
rect 8208 12316 8260 12368
rect 10784 12393 10793 12427
rect 10793 12393 10827 12427
rect 10827 12393 10836 12427
rect 10784 12384 10836 12393
rect 11336 12427 11388 12436
rect 11336 12393 11345 12427
rect 11345 12393 11379 12427
rect 11379 12393 11388 12427
rect 11336 12384 11388 12393
rect 12072 12427 12124 12436
rect 12072 12393 12081 12427
rect 12081 12393 12115 12427
rect 12115 12393 12124 12427
rect 12072 12384 12124 12393
rect 4988 12248 5040 12257
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 5632 12223 5684 12232
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 5632 12180 5684 12189
rect 6184 12180 6236 12232
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 2044 12044 2096 12096
rect 3608 12044 3660 12096
rect 6368 12112 6420 12164
rect 6460 12112 6512 12164
rect 6828 12044 6880 12096
rect 7656 12112 7708 12164
rect 8944 12180 8996 12232
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 8576 12112 8628 12164
rect 8668 12112 8720 12164
rect 9036 12112 9088 12164
rect 9404 12180 9456 12232
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 12348 12316 12400 12368
rect 10692 12291 10744 12300
rect 10692 12257 10701 12291
rect 10701 12257 10735 12291
rect 10735 12257 10744 12291
rect 10692 12248 10744 12257
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 12164 12223 12216 12232
rect 12164 12189 12173 12223
rect 12173 12189 12207 12223
rect 12207 12189 12216 12223
rect 12164 12180 12216 12189
rect 8116 12044 8168 12096
rect 9680 12044 9732 12096
rect 10508 12112 10560 12164
rect 10784 12112 10836 12164
rect 10140 12044 10192 12096
rect 11152 12044 11204 12096
rect 4898 11942 4950 11994
rect 4962 11942 5014 11994
rect 5026 11942 5078 11994
rect 5090 11942 5142 11994
rect 5154 11942 5206 11994
rect 8846 11942 8898 11994
rect 8910 11942 8962 11994
rect 8974 11942 9026 11994
rect 9038 11942 9090 11994
rect 9102 11942 9154 11994
rect 12794 11942 12846 11994
rect 12858 11942 12910 11994
rect 12922 11942 12974 11994
rect 12986 11942 13038 11994
rect 13050 11942 13102 11994
rect 1584 11840 1636 11892
rect 4160 11883 4212 11892
rect 4160 11849 4169 11883
rect 4169 11849 4203 11883
rect 4203 11849 4212 11883
rect 4160 11840 4212 11849
rect 5908 11840 5960 11892
rect 8576 11840 8628 11892
rect 10140 11840 10192 11892
rect 4436 11772 4488 11824
rect 6644 11772 6696 11824
rect 8300 11772 8352 11824
rect 5448 11704 5500 11756
rect 6184 11704 6236 11756
rect 7472 11747 7524 11756
rect 7472 11713 7490 11747
rect 7490 11713 7524 11747
rect 7472 11704 7524 11713
rect 8024 11704 8076 11756
rect 9036 11704 9088 11756
rect 9404 11704 9456 11756
rect 10140 11704 10192 11756
rect 11336 11704 11388 11756
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 12348 11747 12400 11756
rect 2136 11636 2188 11688
rect 2688 11679 2740 11688
rect 2688 11645 2706 11679
rect 2706 11645 2740 11679
rect 2688 11636 2740 11645
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 3516 11679 3568 11688
rect 2780 11636 2832 11645
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 3700 11679 3752 11688
rect 3700 11645 3709 11679
rect 3709 11645 3743 11679
rect 3743 11645 3752 11679
rect 3700 11636 3752 11645
rect 8208 11636 8260 11688
rect 8944 11636 8996 11688
rect 3056 11611 3108 11620
rect 3056 11577 3065 11611
rect 3065 11577 3099 11611
rect 3099 11577 3108 11611
rect 3056 11568 3108 11577
rect 5540 11568 5592 11620
rect 5816 11568 5868 11620
rect 9772 11679 9824 11688
rect 9772 11645 9781 11679
rect 9781 11645 9815 11679
rect 9815 11645 9824 11679
rect 9772 11636 9824 11645
rect 10232 11636 10284 11688
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 2688 11500 2740 11552
rect 7472 11500 7524 11552
rect 8760 11500 8812 11552
rect 8944 11500 8996 11552
rect 9312 11543 9364 11552
rect 9312 11509 9321 11543
rect 9321 11509 9355 11543
rect 9355 11509 9364 11543
rect 9312 11500 9364 11509
rect 11612 11568 11664 11620
rect 11796 11500 11848 11552
rect 2924 11398 2976 11450
rect 2988 11398 3040 11450
rect 3052 11398 3104 11450
rect 3116 11398 3168 11450
rect 3180 11398 3232 11450
rect 6872 11398 6924 11450
rect 6936 11398 6988 11450
rect 7000 11398 7052 11450
rect 7064 11398 7116 11450
rect 7128 11398 7180 11450
rect 10820 11398 10872 11450
rect 10884 11398 10936 11450
rect 10948 11398 11000 11450
rect 11012 11398 11064 11450
rect 11076 11398 11128 11450
rect 14768 11398 14820 11450
rect 14832 11398 14884 11450
rect 14896 11398 14948 11450
rect 14960 11398 15012 11450
rect 15024 11398 15076 11450
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 5632 11339 5684 11348
rect 5632 11305 5641 11339
rect 5641 11305 5675 11339
rect 5675 11305 5684 11339
rect 5632 11296 5684 11305
rect 7380 11296 7432 11348
rect 9864 11296 9916 11348
rect 9956 11296 10008 11348
rect 10324 11296 10376 11348
rect 10784 11296 10836 11348
rect 11612 11339 11664 11348
rect 11612 11305 11621 11339
rect 11621 11305 11655 11339
rect 11655 11305 11664 11339
rect 11612 11296 11664 11305
rect 12624 11296 12676 11348
rect 10048 11228 10100 11280
rect 10508 11228 10560 11280
rect 3424 11092 3476 11144
rect 5448 11160 5500 11212
rect 8024 11203 8076 11212
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 9128 11160 9180 11212
rect 9680 11160 9732 11212
rect 4344 11092 4396 11144
rect 5540 11092 5592 11144
rect 7196 11092 7248 11144
rect 7472 11092 7524 11144
rect 2504 11024 2556 11076
rect 6092 11024 6144 11076
rect 7656 11024 7708 11076
rect 4712 10956 4764 11008
rect 7472 10956 7524 11008
rect 7840 11092 7892 11144
rect 9588 11092 9640 11144
rect 10232 11092 10284 11144
rect 10600 11092 10652 11144
rect 11152 11135 11204 11144
rect 11152 11101 11161 11135
rect 11161 11101 11195 11135
rect 11195 11101 11204 11135
rect 11152 11092 11204 11101
rect 12256 11135 12308 11144
rect 8392 11024 8444 11076
rect 9864 10956 9916 11008
rect 10784 11024 10836 11076
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 12532 11024 12584 11076
rect 12716 11092 12768 11144
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 10876 10956 10928 11008
rect 11244 10999 11296 11008
rect 11244 10965 11253 10999
rect 11253 10965 11287 10999
rect 11287 10965 11296 10999
rect 11244 10956 11296 10965
rect 12072 10999 12124 11008
rect 12072 10965 12081 10999
rect 12081 10965 12115 10999
rect 12115 10965 12124 10999
rect 12072 10956 12124 10965
rect 13360 11024 13412 11076
rect 4898 10854 4950 10906
rect 4962 10854 5014 10906
rect 5026 10854 5078 10906
rect 5090 10854 5142 10906
rect 5154 10854 5206 10906
rect 8846 10854 8898 10906
rect 8910 10854 8962 10906
rect 8974 10854 9026 10906
rect 9038 10854 9090 10906
rect 9102 10854 9154 10906
rect 12794 10854 12846 10906
rect 12858 10854 12910 10906
rect 12922 10854 12974 10906
rect 12986 10854 13038 10906
rect 13050 10854 13102 10906
rect 3516 10752 3568 10804
rect 4068 10684 4120 10736
rect 4252 10684 4304 10736
rect 4896 10684 4948 10736
rect 6552 10752 6604 10804
rect 8116 10752 8168 10804
rect 5908 10684 5960 10736
rect 6368 10684 6420 10736
rect 5356 10616 5408 10668
rect 9312 10684 9364 10736
rect 8300 10616 8352 10668
rect 9680 10752 9732 10804
rect 9772 10752 9824 10804
rect 12164 10752 12216 10804
rect 14096 10752 14148 10804
rect 10324 10659 10376 10668
rect 10324 10625 10333 10659
rect 10333 10625 10367 10659
rect 10367 10625 10376 10659
rect 10324 10616 10376 10625
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 5448 10548 5500 10600
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 10416 10625 10425 10652
rect 10425 10625 10459 10652
rect 10459 10625 10468 10652
rect 10416 10600 10468 10625
rect 10232 10591 10284 10600
rect 3516 10480 3568 10532
rect 4252 10412 4304 10464
rect 6276 10480 6328 10532
rect 7472 10480 7524 10532
rect 10232 10557 10241 10591
rect 10241 10557 10275 10591
rect 10275 10557 10284 10591
rect 10232 10548 10284 10557
rect 10784 10684 10836 10736
rect 11244 10684 11296 10736
rect 12072 10684 12124 10736
rect 12348 10684 12400 10736
rect 13912 10727 13964 10736
rect 12256 10616 12308 10668
rect 12440 10659 12492 10668
rect 12440 10625 12449 10659
rect 12449 10625 12483 10659
rect 12483 10625 12492 10659
rect 12440 10616 12492 10625
rect 12716 10659 12768 10668
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 11428 10480 11480 10532
rect 12072 10548 12124 10600
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 13912 10693 13921 10727
rect 13921 10693 13955 10727
rect 13955 10693 13964 10727
rect 13912 10684 13964 10693
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 14648 10659 14700 10668
rect 13268 10548 13320 10600
rect 14648 10625 14657 10659
rect 14657 10625 14691 10659
rect 14691 10625 14700 10659
rect 14648 10616 14700 10625
rect 12256 10412 12308 10464
rect 12716 10455 12768 10464
rect 12716 10421 12725 10455
rect 12725 10421 12759 10455
rect 12759 10421 12768 10455
rect 12716 10412 12768 10421
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 2924 10310 2976 10362
rect 2988 10310 3040 10362
rect 3052 10310 3104 10362
rect 3116 10310 3168 10362
rect 3180 10310 3232 10362
rect 6872 10310 6924 10362
rect 6936 10310 6988 10362
rect 7000 10310 7052 10362
rect 7064 10310 7116 10362
rect 7128 10310 7180 10362
rect 10820 10310 10872 10362
rect 10884 10310 10936 10362
rect 10948 10310 11000 10362
rect 11012 10310 11064 10362
rect 11076 10310 11128 10362
rect 14768 10310 14820 10362
rect 14832 10310 14884 10362
rect 14896 10310 14948 10362
rect 14960 10310 15012 10362
rect 15024 10310 15076 10362
rect 3700 10208 3752 10260
rect 5540 10072 5592 10124
rect 6368 10208 6420 10260
rect 7288 10208 7340 10260
rect 10600 10208 10652 10260
rect 11520 10208 11572 10260
rect 11888 10208 11940 10260
rect 14096 10251 14148 10260
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 8668 10140 8720 10192
rect 9404 10140 9456 10192
rect 12256 10140 12308 10192
rect 7840 10072 7892 10124
rect 9496 10072 9548 10124
rect 4896 10047 4948 10056
rect 4896 10013 4914 10047
rect 4914 10013 4948 10047
rect 4896 10004 4948 10013
rect 6184 10004 6236 10056
rect 7656 10047 7708 10056
rect 7656 10013 7663 10047
rect 7663 10013 7708 10047
rect 7656 10004 7708 10013
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 8300 10004 8352 10056
rect 9864 10004 9916 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 10784 10004 10836 10056
rect 13268 10072 13320 10124
rect 1768 9979 1820 9988
rect 1768 9945 1777 9979
rect 1777 9945 1811 9979
rect 1811 9945 1820 9979
rect 1768 9936 1820 9945
rect 3332 9936 3384 9988
rect 1584 9868 1636 9920
rect 4436 9936 4488 9988
rect 3608 9868 3660 9920
rect 6276 9936 6328 9988
rect 12072 10004 12124 10056
rect 8392 9868 8444 9920
rect 9680 9911 9732 9920
rect 9680 9877 9689 9911
rect 9689 9877 9723 9911
rect 9723 9877 9732 9911
rect 12624 10004 12676 10056
rect 12716 10004 12768 10056
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 12716 9911 12768 9920
rect 9680 9868 9732 9877
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 4898 9766 4950 9818
rect 4962 9766 5014 9818
rect 5026 9766 5078 9818
rect 5090 9766 5142 9818
rect 5154 9766 5206 9818
rect 8846 9766 8898 9818
rect 8910 9766 8962 9818
rect 8974 9766 9026 9818
rect 9038 9766 9090 9818
rect 9102 9766 9154 9818
rect 12794 9766 12846 9818
rect 12858 9766 12910 9818
rect 12922 9766 12974 9818
rect 12986 9766 13038 9818
rect 13050 9766 13102 9818
rect 1492 9664 1544 9716
rect 4252 9664 4304 9716
rect 3976 9596 4028 9648
rect 5908 9664 5960 9716
rect 7380 9596 7432 9648
rect 8116 9664 8168 9716
rect 9588 9664 9640 9716
rect 4160 9528 4212 9580
rect 7196 9528 7248 9580
rect 3700 9460 3752 9512
rect 3792 9460 3844 9512
rect 4252 9392 4304 9444
rect 3424 9324 3476 9376
rect 4804 9324 4856 9376
rect 6092 9460 6144 9512
rect 6368 9503 6420 9512
rect 6368 9469 6377 9503
rect 6377 9469 6411 9503
rect 6411 9469 6420 9503
rect 6368 9460 6420 9469
rect 7932 9392 7984 9444
rect 8208 9435 8260 9444
rect 8208 9401 8217 9435
rect 8217 9401 8251 9435
rect 8251 9401 8260 9435
rect 8208 9392 8260 9401
rect 8668 9528 8720 9580
rect 9956 9664 10008 9716
rect 10232 9664 10284 9716
rect 12072 9664 12124 9716
rect 12440 9664 12492 9716
rect 13452 9664 13504 9716
rect 9864 9639 9916 9648
rect 9864 9605 9873 9639
rect 9873 9605 9907 9639
rect 9907 9605 9916 9639
rect 9864 9596 9916 9605
rect 11244 9596 11296 9648
rect 8576 9460 8628 9512
rect 9128 9460 9180 9512
rect 9220 9460 9272 9512
rect 10508 9528 10560 9580
rect 13360 9596 13412 9648
rect 12348 9571 12400 9580
rect 10600 9460 10652 9512
rect 12348 9537 12357 9571
rect 12357 9537 12391 9571
rect 12391 9537 12400 9571
rect 12348 9528 12400 9537
rect 12440 9528 12492 9580
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 13268 9571 13320 9580
rect 11612 9460 11664 9512
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 11336 9392 11388 9444
rect 12072 9392 12124 9444
rect 6552 9324 6604 9376
rect 6644 9324 6696 9376
rect 9404 9324 9456 9376
rect 14280 9324 14332 9376
rect 2924 9222 2976 9274
rect 2988 9222 3040 9274
rect 3052 9222 3104 9274
rect 3116 9222 3168 9274
rect 3180 9222 3232 9274
rect 6872 9222 6924 9274
rect 6936 9222 6988 9274
rect 7000 9222 7052 9274
rect 7064 9222 7116 9274
rect 7128 9222 7180 9274
rect 10820 9222 10872 9274
rect 10884 9222 10936 9274
rect 10948 9222 11000 9274
rect 11012 9222 11064 9274
rect 11076 9222 11128 9274
rect 14768 9222 14820 9274
rect 14832 9222 14884 9274
rect 14896 9222 14948 9274
rect 14960 9222 15012 9274
rect 15024 9222 15076 9274
rect 1676 9120 1728 9172
rect 2964 9120 3016 9172
rect 1584 8984 1636 9036
rect 4252 9120 4304 9172
rect 6460 9120 6512 9172
rect 6552 9120 6604 9172
rect 7932 9120 7984 9172
rect 9772 9120 9824 9172
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 10508 9120 10560 9172
rect 4528 8984 4580 9036
rect 4620 8984 4672 9036
rect 7288 9052 7340 9104
rect 7656 9052 7708 9104
rect 6276 9027 6328 9036
rect 6276 8993 6285 9027
rect 6285 8993 6319 9027
rect 6319 8993 6328 9027
rect 6276 8984 6328 8993
rect 9588 9052 9640 9104
rect 2320 8848 2372 8900
rect 3516 8916 3568 8968
rect 3424 8848 3476 8900
rect 1676 8780 1728 8832
rect 2964 8780 3016 8832
rect 5448 8848 5500 8900
rect 6092 8916 6144 8968
rect 7472 8916 7524 8968
rect 6276 8848 6328 8900
rect 5908 8780 5960 8832
rect 7472 8780 7524 8832
rect 7748 8780 7800 8832
rect 8208 8916 8260 8968
rect 8484 8984 8536 9036
rect 8576 8916 8628 8968
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9496 8959 9548 8968
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 9496 8916 9548 8925
rect 9036 8848 9088 8900
rect 10600 9052 10652 9104
rect 11152 9120 11204 9172
rect 12624 9052 12676 9104
rect 11060 8984 11112 9036
rect 10600 8916 10652 8968
rect 12072 8984 12124 9036
rect 10416 8848 10468 8900
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11980 8959 12032 8968
rect 11336 8916 11388 8925
rect 11980 8925 11989 8959
rect 11989 8925 12023 8959
rect 12023 8925 12032 8959
rect 11980 8916 12032 8925
rect 12624 8959 12676 8968
rect 11152 8848 11204 8900
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 8024 8780 8076 8832
rect 8484 8780 8536 8832
rect 9312 8780 9364 8832
rect 10048 8780 10100 8832
rect 10508 8780 10560 8832
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 11244 8823 11296 8832
rect 11244 8789 11253 8823
rect 11253 8789 11287 8823
rect 11287 8789 11296 8823
rect 11244 8780 11296 8789
rect 11704 8780 11756 8832
rect 4898 8678 4950 8730
rect 4962 8678 5014 8730
rect 5026 8678 5078 8730
rect 5090 8678 5142 8730
rect 5154 8678 5206 8730
rect 8846 8678 8898 8730
rect 8910 8678 8962 8730
rect 8974 8678 9026 8730
rect 9038 8678 9090 8730
rect 9102 8678 9154 8730
rect 12794 8678 12846 8730
rect 12858 8678 12910 8730
rect 12922 8678 12974 8730
rect 12986 8678 13038 8730
rect 13050 8678 13102 8730
rect 6828 8576 6880 8628
rect 7564 8576 7616 8628
rect 5264 8508 5316 8560
rect 9496 8576 9548 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 3516 8440 3568 8492
rect 8484 8508 8536 8560
rect 9036 8508 9088 8560
rect 10508 8576 10560 8628
rect 11796 8576 11848 8628
rect 12164 8619 12216 8628
rect 12164 8585 12173 8619
rect 12173 8585 12207 8619
rect 12207 8585 12216 8619
rect 12164 8576 12216 8585
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 4712 8372 4764 8424
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 7104 8440 7156 8492
rect 8024 8440 8076 8492
rect 6552 8415 6604 8424
rect 5080 8304 5132 8356
rect 6000 8304 6052 8356
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 7564 8347 7616 8356
rect 7564 8313 7573 8347
rect 7573 8313 7607 8347
rect 7607 8313 7616 8347
rect 7564 8304 7616 8313
rect 8024 8304 8076 8356
rect 8668 8440 8720 8492
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 9496 8440 9548 8492
rect 9772 8440 9824 8492
rect 4712 8236 4764 8288
rect 6552 8236 6604 8288
rect 10416 8372 10468 8424
rect 10968 8508 11020 8560
rect 11428 8508 11480 8560
rect 10692 8440 10744 8492
rect 10876 8440 10928 8492
rect 11612 8440 11664 8492
rect 12348 8483 12400 8492
rect 12348 8449 12357 8483
rect 12357 8449 12391 8483
rect 12391 8449 12400 8483
rect 12348 8440 12400 8449
rect 8668 8347 8720 8356
rect 8668 8313 8677 8347
rect 8677 8313 8711 8347
rect 8711 8313 8720 8347
rect 8668 8304 8720 8313
rect 8760 8304 8812 8356
rect 9496 8236 9548 8288
rect 10508 8304 10560 8356
rect 14648 8372 14700 8424
rect 12440 8304 12492 8356
rect 10784 8236 10836 8288
rect 11060 8236 11112 8288
rect 11244 8236 11296 8288
rect 2924 8134 2976 8186
rect 2988 8134 3040 8186
rect 3052 8134 3104 8186
rect 3116 8134 3168 8186
rect 3180 8134 3232 8186
rect 6872 8134 6924 8186
rect 6936 8134 6988 8186
rect 7000 8134 7052 8186
rect 7064 8134 7116 8186
rect 7128 8134 7180 8186
rect 10820 8134 10872 8186
rect 10884 8134 10936 8186
rect 10948 8134 11000 8186
rect 11012 8134 11064 8186
rect 11076 8134 11128 8186
rect 14768 8134 14820 8186
rect 14832 8134 14884 8186
rect 14896 8134 14948 8186
rect 14960 8134 15012 8186
rect 15024 8134 15076 8186
rect 4252 8032 4304 8084
rect 4712 8032 4764 8084
rect 3240 7896 3292 7948
rect 6000 7896 6052 7948
rect 2780 7828 2832 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 5632 7828 5684 7880
rect 6276 7828 6328 7880
rect 6368 7828 6420 7880
rect 7104 7964 7156 8016
rect 7656 8032 7708 8084
rect 7840 8032 7892 8084
rect 8300 8075 8352 8084
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 9404 8032 9456 8084
rect 11888 8075 11940 8084
rect 11888 8041 11897 8075
rect 11897 8041 11931 8075
rect 11931 8041 11940 8075
rect 11888 8032 11940 8041
rect 8116 7964 8168 8016
rect 8484 7964 8536 8016
rect 9220 7964 9272 8016
rect 13176 7964 13228 8016
rect 6828 7896 6880 7948
rect 7840 7896 7892 7948
rect 7104 7828 7156 7880
rect 7932 7828 7984 7880
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 10600 7828 10652 7880
rect 10968 7828 11020 7880
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 12440 7896 12492 7948
rect 12624 7896 12676 7948
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 1676 7803 1728 7812
rect 1676 7769 1685 7803
rect 1685 7769 1719 7803
rect 1719 7769 1728 7803
rect 1676 7760 1728 7769
rect 4068 7803 4120 7812
rect 4068 7769 4077 7803
rect 4077 7769 4111 7803
rect 4111 7769 4120 7803
rect 4068 7760 4120 7769
rect 5448 7760 5500 7812
rect 9404 7803 9456 7812
rect 9404 7769 9413 7803
rect 9413 7769 9447 7803
rect 9447 7769 9456 7803
rect 9404 7760 9456 7769
rect 1584 7692 1636 7744
rect 2688 7692 2740 7744
rect 3516 7692 3568 7744
rect 5080 7692 5132 7744
rect 5908 7692 5960 7744
rect 6368 7735 6420 7744
rect 6368 7701 6377 7735
rect 6377 7701 6411 7735
rect 6411 7701 6420 7735
rect 6368 7692 6420 7701
rect 7012 7692 7064 7744
rect 7288 7692 7340 7744
rect 8300 7692 8352 7744
rect 9864 7692 9916 7744
rect 11060 7692 11112 7744
rect 11244 7692 11296 7744
rect 4898 7590 4950 7642
rect 4962 7590 5014 7642
rect 5026 7590 5078 7642
rect 5090 7590 5142 7642
rect 5154 7590 5206 7642
rect 8846 7590 8898 7642
rect 8910 7590 8962 7642
rect 8974 7590 9026 7642
rect 9038 7590 9090 7642
rect 9102 7590 9154 7642
rect 12794 7590 12846 7642
rect 12858 7590 12910 7642
rect 12922 7590 12974 7642
rect 12986 7590 13038 7642
rect 13050 7590 13102 7642
rect 3516 7488 3568 7540
rect 3240 7420 3292 7472
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 3056 7352 3108 7404
rect 3884 7420 3936 7472
rect 3516 7352 3568 7404
rect 3976 7395 4028 7404
rect 3976 7361 4010 7395
rect 4010 7361 4028 7395
rect 3976 7352 4028 7361
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 2412 7284 2464 7336
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 5908 7352 5960 7404
rect 7196 7488 7248 7540
rect 7288 7488 7340 7540
rect 8760 7531 8812 7540
rect 5724 7284 5776 7336
rect 6736 7395 6788 7404
rect 6736 7361 6769 7395
rect 6769 7361 6788 7395
rect 7012 7420 7064 7472
rect 8392 7463 8444 7472
rect 8392 7429 8401 7463
rect 8401 7429 8435 7463
rect 8435 7429 8444 7463
rect 8392 7420 8444 7429
rect 8760 7497 8769 7531
rect 8769 7497 8803 7531
rect 8803 7497 8812 7531
rect 8760 7488 8812 7497
rect 6736 7352 6788 7361
rect 7288 7352 7340 7404
rect 7656 7352 7708 7404
rect 8760 7352 8812 7404
rect 8944 7420 8996 7472
rect 10232 7488 10284 7540
rect 10416 7488 10468 7540
rect 9680 7420 9732 7472
rect 6460 7284 6512 7336
rect 7472 7327 7524 7336
rect 7472 7293 7481 7327
rect 7481 7293 7515 7327
rect 7515 7293 7524 7327
rect 7472 7284 7524 7293
rect 8944 7284 8996 7336
rect 9772 7352 9824 7404
rect 11612 7420 11664 7472
rect 10048 7395 10100 7404
rect 10048 7361 10057 7395
rect 10057 7361 10091 7395
rect 10091 7361 10100 7395
rect 10508 7395 10560 7404
rect 10048 7352 10100 7361
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 10600 7352 10652 7404
rect 4712 7216 4764 7268
rect 9128 7216 9180 7268
rect 12348 7284 12400 7336
rect 12256 7216 12308 7268
rect 2136 7148 2188 7200
rect 3056 7148 3108 7200
rect 3516 7148 3568 7200
rect 4988 7148 5040 7200
rect 9404 7148 9456 7200
rect 2924 7046 2976 7098
rect 2988 7046 3040 7098
rect 3052 7046 3104 7098
rect 3116 7046 3168 7098
rect 3180 7046 3232 7098
rect 6872 7046 6924 7098
rect 6936 7046 6988 7098
rect 7000 7046 7052 7098
rect 7064 7046 7116 7098
rect 7128 7046 7180 7098
rect 10820 7046 10872 7098
rect 10884 7046 10936 7098
rect 10948 7046 11000 7098
rect 11012 7046 11064 7098
rect 11076 7046 11128 7098
rect 14768 7046 14820 7098
rect 14832 7046 14884 7098
rect 14896 7046 14948 7098
rect 14960 7046 15012 7098
rect 15024 7046 15076 7098
rect 1492 6944 1544 6996
rect 4068 6944 4120 6996
rect 5172 6987 5224 6996
rect 5172 6953 5181 6987
rect 5181 6953 5215 6987
rect 5215 6953 5224 6987
rect 5172 6944 5224 6953
rect 5632 6987 5684 6996
rect 5632 6953 5641 6987
rect 5641 6953 5675 6987
rect 5675 6953 5684 6987
rect 5632 6944 5684 6953
rect 2872 6876 2924 6928
rect 3884 6876 3936 6928
rect 4160 6876 4212 6928
rect 5540 6876 5592 6928
rect 6000 6944 6052 6996
rect 6092 6987 6144 6996
rect 6092 6953 6101 6987
rect 6101 6953 6135 6987
rect 6135 6953 6144 6987
rect 6092 6944 6144 6953
rect 6368 6944 6420 6996
rect 6828 6944 6880 6996
rect 7012 6944 7064 6996
rect 8760 6944 8812 6996
rect 9036 6987 9088 6996
rect 9036 6953 9045 6987
rect 9045 6953 9079 6987
rect 9079 6953 9088 6987
rect 9036 6944 9088 6953
rect 9588 6987 9640 6996
rect 9588 6953 9597 6987
rect 9597 6953 9631 6987
rect 9631 6953 9640 6987
rect 9588 6944 9640 6953
rect 6736 6876 6788 6928
rect 9312 6876 9364 6928
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 3148 6808 3200 6860
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 4436 6808 4488 6860
rect 7472 6808 7524 6860
rect 7564 6851 7616 6860
rect 7564 6817 7573 6851
rect 7573 6817 7607 6851
rect 7607 6817 7616 6851
rect 7564 6808 7616 6817
rect 4252 6740 4304 6792
rect 6552 6740 6604 6792
rect 6920 6740 6972 6792
rect 3792 6604 3844 6656
rect 4068 6604 4120 6656
rect 4436 6604 4488 6656
rect 4988 6604 5040 6656
rect 5816 6672 5868 6724
rect 6736 6672 6788 6724
rect 7012 6672 7064 6724
rect 7748 6740 7800 6792
rect 7932 6740 7984 6792
rect 8668 6808 8720 6860
rect 8116 6672 8168 6724
rect 8392 6740 8444 6792
rect 10140 6808 10192 6860
rect 9220 6740 9272 6792
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 11428 6740 11480 6792
rect 6000 6604 6052 6656
rect 6276 6604 6328 6656
rect 6460 6604 6512 6656
rect 9956 6604 10008 6656
rect 4898 6502 4950 6554
rect 4962 6502 5014 6554
rect 5026 6502 5078 6554
rect 5090 6502 5142 6554
rect 5154 6502 5206 6554
rect 8846 6502 8898 6554
rect 8910 6502 8962 6554
rect 8974 6502 9026 6554
rect 9038 6502 9090 6554
rect 9102 6502 9154 6554
rect 12794 6502 12846 6554
rect 12858 6502 12910 6554
rect 12922 6502 12974 6554
rect 12986 6502 13038 6554
rect 13050 6502 13102 6554
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 2780 6400 2832 6409
rect 1860 6332 1912 6384
rect 2412 6332 2464 6384
rect 4988 6400 5040 6452
rect 5356 6400 5408 6452
rect 5816 6400 5868 6452
rect 6368 6443 6420 6452
rect 6368 6409 6377 6443
rect 6377 6409 6411 6443
rect 6411 6409 6420 6443
rect 6368 6400 6420 6409
rect 6828 6400 6880 6452
rect 4436 6332 4488 6384
rect 4712 6375 4764 6384
rect 1492 6264 1544 6316
rect 1952 6264 2004 6316
rect 3148 6264 3200 6316
rect 4252 6264 4304 6316
rect 4712 6341 4721 6375
rect 4721 6341 4755 6375
rect 4755 6341 4764 6375
rect 4712 6332 4764 6341
rect 3516 6196 3568 6248
rect 4344 6196 4396 6248
rect 3792 6128 3844 6180
rect 3516 6060 3568 6112
rect 5080 6264 5132 6316
rect 5356 6264 5408 6316
rect 5632 6264 5684 6316
rect 6092 6332 6144 6384
rect 6276 6332 6328 6384
rect 10692 6400 10744 6452
rect 4988 6196 5040 6248
rect 6092 6196 6144 6248
rect 7196 6264 7248 6316
rect 7748 6332 7800 6384
rect 9220 6332 9272 6384
rect 10048 6332 10100 6384
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 8576 6264 8628 6316
rect 8668 6196 8720 6248
rect 9588 6196 9640 6248
rect 5080 6128 5132 6180
rect 6000 6128 6052 6180
rect 7840 6128 7892 6180
rect 8760 6171 8812 6180
rect 8760 6137 8769 6171
rect 8769 6137 8803 6171
rect 8803 6137 8812 6171
rect 8760 6128 8812 6137
rect 7196 6060 7248 6112
rect 7481 6103 7533 6112
rect 7481 6069 7490 6103
rect 7490 6069 7524 6103
rect 7524 6069 7533 6103
rect 7481 6060 7533 6069
rect 8116 6060 8168 6112
rect 11152 6060 11204 6112
rect 2924 5958 2976 6010
rect 2988 5958 3040 6010
rect 3052 5958 3104 6010
rect 3116 5958 3168 6010
rect 3180 5958 3232 6010
rect 6872 5958 6924 6010
rect 6936 5958 6988 6010
rect 7000 5958 7052 6010
rect 7064 5958 7116 6010
rect 7128 5958 7180 6010
rect 10820 5958 10872 6010
rect 10884 5958 10936 6010
rect 10948 5958 11000 6010
rect 11012 5958 11064 6010
rect 11076 5958 11128 6010
rect 14768 5958 14820 6010
rect 14832 5958 14884 6010
rect 14896 5958 14948 6010
rect 14960 5958 15012 6010
rect 15024 5958 15076 6010
rect 4528 5856 4580 5908
rect 6552 5856 6604 5908
rect 3792 5788 3844 5840
rect 7564 5788 7616 5840
rect 1768 5720 1820 5772
rect 2596 5652 2648 5704
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4528 5720 4580 5772
rect 5632 5763 5684 5772
rect 3976 5584 4028 5636
rect 4252 5584 4304 5636
rect 5356 5652 5408 5704
rect 5632 5729 5641 5763
rect 5641 5729 5675 5763
rect 5675 5729 5684 5763
rect 5632 5720 5684 5729
rect 7288 5720 7340 5772
rect 6736 5652 6788 5704
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7380 5652 7432 5704
rect 8484 5720 8536 5772
rect 9680 5720 9732 5772
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 7840 5652 7892 5704
rect 10508 5652 10560 5704
rect 6092 5627 6144 5636
rect 6092 5593 6101 5627
rect 6101 5593 6135 5627
rect 6135 5593 6144 5627
rect 6092 5584 6144 5593
rect 2596 5516 2648 5568
rect 10600 5584 10652 5636
rect 6276 5559 6328 5568
rect 6276 5525 6301 5559
rect 6301 5525 6328 5559
rect 6276 5516 6328 5525
rect 7104 5516 7156 5568
rect 7380 5516 7432 5568
rect 8024 5516 8076 5568
rect 8484 5516 8536 5568
rect 4898 5414 4950 5466
rect 4962 5414 5014 5466
rect 5026 5414 5078 5466
rect 5090 5414 5142 5466
rect 5154 5414 5206 5466
rect 8846 5414 8898 5466
rect 8910 5414 8962 5466
rect 8974 5414 9026 5466
rect 9038 5414 9090 5466
rect 9102 5414 9154 5466
rect 12794 5414 12846 5466
rect 12858 5414 12910 5466
rect 12922 5414 12974 5466
rect 12986 5414 13038 5466
rect 13050 5414 13102 5466
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 5356 5312 5408 5364
rect 5540 5312 5592 5364
rect 6276 5312 6328 5364
rect 6460 5355 6512 5364
rect 6460 5321 6469 5355
rect 6469 5321 6503 5355
rect 6503 5321 6512 5355
rect 6460 5312 6512 5321
rect 6920 5312 6972 5364
rect 7196 5312 7248 5364
rect 11980 5312 12032 5364
rect 3516 5244 3568 5296
rect 2504 5176 2556 5228
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 3976 5176 4028 5228
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 4252 5176 4304 5185
rect 6092 5244 6144 5296
rect 5540 5176 5592 5228
rect 5724 5176 5776 5228
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 8484 5244 8536 5296
rect 6368 5176 6420 5185
rect 6736 5176 6788 5228
rect 7104 5176 7156 5228
rect 11520 5176 11572 5228
rect 2596 5151 2648 5160
rect 2596 5117 2605 5151
rect 2605 5117 2639 5151
rect 2639 5117 2648 5151
rect 2596 5108 2648 5117
rect 4528 5108 4580 5160
rect 5908 5108 5960 5160
rect 6000 5108 6052 5160
rect 8116 5108 8168 5160
rect 4068 5040 4120 5092
rect 6736 5040 6788 5092
rect 7288 5040 7340 5092
rect 11796 5040 11848 5092
rect 4712 4972 4764 5024
rect 4804 4972 4856 5024
rect 5356 4972 5408 5024
rect 6184 4972 6236 5024
rect 6368 4972 6420 5024
rect 8208 4972 8260 5024
rect 2924 4870 2976 4922
rect 2988 4870 3040 4922
rect 3052 4870 3104 4922
rect 3116 4870 3168 4922
rect 3180 4870 3232 4922
rect 6872 4870 6924 4922
rect 6936 4870 6988 4922
rect 7000 4870 7052 4922
rect 7064 4870 7116 4922
rect 7128 4870 7180 4922
rect 10820 4870 10872 4922
rect 10884 4870 10936 4922
rect 10948 4870 11000 4922
rect 11012 4870 11064 4922
rect 11076 4870 11128 4922
rect 14768 4870 14820 4922
rect 14832 4870 14884 4922
rect 14896 4870 14948 4922
rect 14960 4870 15012 4922
rect 15024 4870 15076 4922
rect 3056 4811 3108 4820
rect 3056 4777 3065 4811
rect 3065 4777 3099 4811
rect 3099 4777 3108 4811
rect 3056 4768 3108 4777
rect 4068 4768 4120 4820
rect 4528 4768 4580 4820
rect 5540 4700 5592 4752
rect 5816 4768 5868 4820
rect 6184 4768 6236 4820
rect 6552 4700 6604 4752
rect 6736 4768 6788 4820
rect 9496 4700 9548 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 1676 4675 1728 4684
rect 1676 4641 1685 4675
rect 1685 4641 1719 4675
rect 1719 4641 1728 4675
rect 1676 4632 1728 4641
rect 2688 4564 2740 4616
rect 4436 4632 4488 4684
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4988 4632 5040 4684
rect 7196 4632 7248 4684
rect 4068 4564 4120 4573
rect 4620 4564 4672 4616
rect 2228 4428 2280 4480
rect 4344 4496 4396 4548
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 4988 4496 5040 4548
rect 4160 4428 4212 4480
rect 5356 4428 5408 4480
rect 12440 4496 12492 4548
rect 9864 4428 9916 4480
rect 4898 4326 4950 4378
rect 4962 4326 5014 4378
rect 5026 4326 5078 4378
rect 5090 4326 5142 4378
rect 5154 4326 5206 4378
rect 8846 4326 8898 4378
rect 8910 4326 8962 4378
rect 8974 4326 9026 4378
rect 9038 4326 9090 4378
rect 9102 4326 9154 4378
rect 12794 4326 12846 4378
rect 12858 4326 12910 4378
rect 12922 4326 12974 4378
rect 12986 4326 13038 4378
rect 13050 4326 13102 4378
rect 2872 4224 2924 4276
rect 2964 4224 3016 4276
rect 7748 4224 7800 4276
rect 3608 4199 3660 4208
rect 3608 4165 3617 4199
rect 3617 4165 3651 4199
rect 3651 4165 3660 4199
rect 3608 4156 3660 4165
rect 4252 4156 4304 4208
rect 1768 4088 1820 4140
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 4528 4156 4580 4208
rect 6000 4156 6052 4208
rect 4620 4131 4672 4140
rect 1400 4063 1452 4072
rect 1400 4029 1409 4063
rect 1409 4029 1443 4063
rect 1443 4029 1452 4063
rect 1400 4020 1452 4029
rect 2504 4020 2556 4072
rect 2964 4020 3016 4072
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 5080 4131 5132 4140
rect 5080 4097 5089 4131
rect 5089 4097 5123 4131
rect 5123 4097 5132 4131
rect 5080 4088 5132 4097
rect 3976 4063 4028 4072
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 6184 4088 6236 4140
rect 3884 3952 3936 4004
rect 5264 3952 5316 4004
rect 4344 3884 4396 3936
rect 7380 3884 7432 3936
rect 2924 3782 2976 3834
rect 2988 3782 3040 3834
rect 3052 3782 3104 3834
rect 3116 3782 3168 3834
rect 3180 3782 3232 3834
rect 6872 3782 6924 3834
rect 6936 3782 6988 3834
rect 7000 3782 7052 3834
rect 7064 3782 7116 3834
rect 7128 3782 7180 3834
rect 10820 3782 10872 3834
rect 10884 3782 10936 3834
rect 10948 3782 11000 3834
rect 11012 3782 11064 3834
rect 11076 3782 11128 3834
rect 14768 3782 14820 3834
rect 14832 3782 14884 3834
rect 14896 3782 14948 3834
rect 14960 3782 15012 3834
rect 15024 3782 15076 3834
rect 2320 3680 2372 3732
rect 4344 3680 4396 3732
rect 11244 3680 11296 3732
rect 2044 3544 2096 3596
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 2688 3612 2740 3664
rect 2228 3519 2280 3528
rect 2228 3485 2237 3519
rect 2237 3485 2271 3519
rect 2271 3485 2280 3519
rect 2228 3476 2280 3485
rect 3700 3612 3752 3664
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 3056 3476 3108 3528
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 3884 3476 3936 3528
rect 5080 3544 5132 3596
rect 8300 3476 8352 3528
rect 2136 3340 2188 3392
rect 11336 3408 11388 3460
rect 4068 3340 4120 3392
rect 4898 3238 4950 3290
rect 4962 3238 5014 3290
rect 5026 3238 5078 3290
rect 5090 3238 5142 3290
rect 5154 3238 5206 3290
rect 8846 3238 8898 3290
rect 8910 3238 8962 3290
rect 8974 3238 9026 3290
rect 9038 3238 9090 3290
rect 9102 3238 9154 3290
rect 12794 3238 12846 3290
rect 12858 3238 12910 3290
rect 12922 3238 12974 3290
rect 12986 3238 13038 3290
rect 13050 3238 13102 3290
rect 2412 3179 2464 3188
rect 2412 3145 2421 3179
rect 2421 3145 2455 3179
rect 2455 3145 2464 3179
rect 2412 3136 2464 3145
rect 3332 3136 3384 3188
rect 1860 3068 1912 3120
rect 3148 3068 3200 3120
rect 1584 3000 1636 3052
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 2504 3000 2556 3052
rect 7932 3000 7984 3052
rect 8392 2932 8444 2984
rect 3148 2864 3200 2916
rect 9772 2796 9824 2848
rect 2924 2694 2976 2746
rect 2988 2694 3040 2746
rect 3052 2694 3104 2746
rect 3116 2694 3168 2746
rect 3180 2694 3232 2746
rect 6872 2694 6924 2746
rect 6936 2694 6988 2746
rect 7000 2694 7052 2746
rect 7064 2694 7116 2746
rect 7128 2694 7180 2746
rect 10820 2694 10872 2746
rect 10884 2694 10936 2746
rect 10948 2694 11000 2746
rect 11012 2694 11064 2746
rect 11076 2694 11128 2746
rect 14768 2694 14820 2746
rect 14832 2694 14884 2746
rect 14896 2694 14948 2746
rect 14960 2694 15012 2746
rect 15024 2694 15076 2746
rect 1952 2592 2004 2644
rect 2688 2524 2740 2576
rect 2044 2456 2096 2508
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 5724 2388 5776 2440
rect 4898 2150 4950 2202
rect 4962 2150 5014 2202
rect 5026 2150 5078 2202
rect 5090 2150 5142 2202
rect 5154 2150 5206 2202
rect 8846 2150 8898 2202
rect 8910 2150 8962 2202
rect 8974 2150 9026 2202
rect 9038 2150 9090 2202
rect 9102 2150 9154 2202
rect 12794 2150 12846 2202
rect 12858 2150 12910 2202
rect 12922 2150 12974 2202
rect 12986 2150 13038 2202
rect 13050 2150 13102 2202
rect 3608 2048 3660 2100
rect 3424 1980 3476 2032
rect 2044 1955 2096 1964
rect 2044 1921 2053 1955
rect 2053 1921 2087 1955
rect 2087 1921 2096 1955
rect 2044 1912 2096 1921
rect 2688 1912 2740 1964
rect 2780 1844 2832 1896
rect 2924 1606 2976 1658
rect 2988 1606 3040 1658
rect 3052 1606 3104 1658
rect 3116 1606 3168 1658
rect 3180 1606 3232 1658
rect 6872 1606 6924 1658
rect 6936 1606 6988 1658
rect 7000 1606 7052 1658
rect 7064 1606 7116 1658
rect 7128 1606 7180 1658
rect 10820 1606 10872 1658
rect 10884 1606 10936 1658
rect 10948 1606 11000 1658
rect 11012 1606 11064 1658
rect 11076 1606 11128 1658
rect 14768 1606 14820 1658
rect 14832 1606 14884 1658
rect 14896 1606 14948 1658
rect 14960 1606 15012 1658
rect 15024 1606 15076 1658
rect 1400 1343 1452 1352
rect 1400 1309 1409 1343
rect 1409 1309 1443 1343
rect 1443 1309 1452 1343
rect 1400 1300 1452 1309
rect 1492 1164 1544 1216
rect 4898 1062 4950 1114
rect 4962 1062 5014 1114
rect 5026 1062 5078 1114
rect 5090 1062 5142 1114
rect 5154 1062 5206 1114
rect 8846 1062 8898 1114
rect 8910 1062 8962 1114
rect 8974 1062 9026 1114
rect 9038 1062 9090 1114
rect 9102 1062 9154 1114
rect 12794 1062 12846 1114
rect 12858 1062 12910 1114
rect 12922 1062 12974 1114
rect 12986 1062 13038 1114
rect 13050 1062 13102 1114
<< metal2 >>
rect 2778 23216 2834 23225
rect 2778 23151 2834 23160
rect 1490 21720 1546 21729
rect 1490 21655 1546 21664
rect 1504 18970 1532 21655
rect 2792 20602 2820 23151
rect 4898 22876 5206 22885
rect 4898 22874 4904 22876
rect 4960 22874 4984 22876
rect 5040 22874 5064 22876
rect 5120 22874 5144 22876
rect 5200 22874 5206 22876
rect 4960 22822 4962 22874
rect 5142 22822 5144 22874
rect 4898 22820 4904 22822
rect 4960 22820 4984 22822
rect 5040 22820 5064 22822
rect 5120 22820 5144 22822
rect 5200 22820 5206 22822
rect 4898 22811 5206 22820
rect 8846 22876 9154 22885
rect 8846 22874 8852 22876
rect 8908 22874 8932 22876
rect 8988 22874 9012 22876
rect 9068 22874 9092 22876
rect 9148 22874 9154 22876
rect 8908 22822 8910 22874
rect 9090 22822 9092 22874
rect 8846 22820 8852 22822
rect 8908 22820 8932 22822
rect 8988 22820 9012 22822
rect 9068 22820 9092 22822
rect 9148 22820 9154 22822
rect 8846 22811 9154 22820
rect 12794 22876 13102 22885
rect 12794 22874 12800 22876
rect 12856 22874 12880 22876
rect 12936 22874 12960 22876
rect 13016 22874 13040 22876
rect 13096 22874 13102 22876
rect 12856 22822 12858 22874
rect 13038 22822 13040 22874
rect 12794 22820 12800 22822
rect 12856 22820 12880 22822
rect 12936 22820 12960 22822
rect 13016 22820 13040 22822
rect 13096 22820 13102 22822
rect 12794 22811 13102 22820
rect 2924 22332 3232 22341
rect 2924 22330 2930 22332
rect 2986 22330 3010 22332
rect 3066 22330 3090 22332
rect 3146 22330 3170 22332
rect 3226 22330 3232 22332
rect 2986 22278 2988 22330
rect 3168 22278 3170 22330
rect 2924 22276 2930 22278
rect 2986 22276 3010 22278
rect 3066 22276 3090 22278
rect 3146 22276 3170 22278
rect 3226 22276 3232 22278
rect 2924 22267 3232 22276
rect 6872 22332 7180 22341
rect 6872 22330 6878 22332
rect 6934 22330 6958 22332
rect 7014 22330 7038 22332
rect 7094 22330 7118 22332
rect 7174 22330 7180 22332
rect 6934 22278 6936 22330
rect 7116 22278 7118 22330
rect 6872 22276 6878 22278
rect 6934 22276 6958 22278
rect 7014 22276 7038 22278
rect 7094 22276 7118 22278
rect 7174 22276 7180 22278
rect 6872 22267 7180 22276
rect 10820 22332 11128 22341
rect 10820 22330 10826 22332
rect 10882 22330 10906 22332
rect 10962 22330 10986 22332
rect 11042 22330 11066 22332
rect 11122 22330 11128 22332
rect 10882 22278 10884 22330
rect 11064 22278 11066 22330
rect 10820 22276 10826 22278
rect 10882 22276 10906 22278
rect 10962 22276 10986 22278
rect 11042 22276 11066 22278
rect 11122 22276 11128 22278
rect 10820 22267 11128 22276
rect 14768 22332 15076 22341
rect 14768 22330 14774 22332
rect 14830 22330 14854 22332
rect 14910 22330 14934 22332
rect 14990 22330 15014 22332
rect 15070 22330 15076 22332
rect 14830 22278 14832 22330
rect 15012 22278 15014 22330
rect 14768 22276 14774 22278
rect 14830 22276 14854 22278
rect 14910 22276 14934 22278
rect 14990 22276 15014 22278
rect 15070 22276 15076 22278
rect 14768 22267 15076 22276
rect 4898 21788 5206 21797
rect 4898 21786 4904 21788
rect 4960 21786 4984 21788
rect 5040 21786 5064 21788
rect 5120 21786 5144 21788
rect 5200 21786 5206 21788
rect 4960 21734 4962 21786
rect 5142 21734 5144 21786
rect 4898 21732 4904 21734
rect 4960 21732 4984 21734
rect 5040 21732 5064 21734
rect 5120 21732 5144 21734
rect 5200 21732 5206 21734
rect 4898 21723 5206 21732
rect 8846 21788 9154 21797
rect 8846 21786 8852 21788
rect 8908 21786 8932 21788
rect 8988 21786 9012 21788
rect 9068 21786 9092 21788
rect 9148 21786 9154 21788
rect 8908 21734 8910 21786
rect 9090 21734 9092 21786
rect 8846 21732 8852 21734
rect 8908 21732 8932 21734
rect 8988 21732 9012 21734
rect 9068 21732 9092 21734
rect 9148 21732 9154 21734
rect 8846 21723 9154 21732
rect 12794 21788 13102 21797
rect 12794 21786 12800 21788
rect 12856 21786 12880 21788
rect 12936 21786 12960 21788
rect 13016 21786 13040 21788
rect 13096 21786 13102 21788
rect 12856 21734 12858 21786
rect 13038 21734 13040 21786
rect 12794 21732 12800 21734
rect 12856 21732 12880 21734
rect 12936 21732 12960 21734
rect 13016 21732 13040 21734
rect 13096 21732 13102 21734
rect 12794 21723 13102 21732
rect 2924 21244 3232 21253
rect 2924 21242 2930 21244
rect 2986 21242 3010 21244
rect 3066 21242 3090 21244
rect 3146 21242 3170 21244
rect 3226 21242 3232 21244
rect 2986 21190 2988 21242
rect 3168 21190 3170 21242
rect 2924 21188 2930 21190
rect 2986 21188 3010 21190
rect 3066 21188 3090 21190
rect 3146 21188 3170 21190
rect 3226 21188 3232 21190
rect 2924 21179 3232 21188
rect 6872 21244 7180 21253
rect 6872 21242 6878 21244
rect 6934 21242 6958 21244
rect 7014 21242 7038 21244
rect 7094 21242 7118 21244
rect 7174 21242 7180 21244
rect 6934 21190 6936 21242
rect 7116 21190 7118 21242
rect 6872 21188 6878 21190
rect 6934 21188 6958 21190
rect 7014 21188 7038 21190
rect 7094 21188 7118 21190
rect 7174 21188 7180 21190
rect 6872 21179 7180 21188
rect 10820 21244 11128 21253
rect 10820 21242 10826 21244
rect 10882 21242 10906 21244
rect 10962 21242 10986 21244
rect 11042 21242 11066 21244
rect 11122 21242 11128 21244
rect 10882 21190 10884 21242
rect 11064 21190 11066 21242
rect 10820 21188 10826 21190
rect 10882 21188 10906 21190
rect 10962 21188 10986 21190
rect 11042 21188 11066 21190
rect 11122 21188 11128 21190
rect 10820 21179 11128 21188
rect 14768 21244 15076 21253
rect 14768 21242 14774 21244
rect 14830 21242 14854 21244
rect 14910 21242 14934 21244
rect 14990 21242 15014 21244
rect 15070 21242 15076 21244
rect 14830 21190 14832 21242
rect 15012 21190 15014 21242
rect 14768 21188 14774 21190
rect 14830 21188 14854 21190
rect 14910 21188 14934 21190
rect 14990 21188 15014 21190
rect 15070 21188 15076 21190
rect 14768 21179 15076 21188
rect 4898 20700 5206 20709
rect 4898 20698 4904 20700
rect 4960 20698 4984 20700
rect 5040 20698 5064 20700
rect 5120 20698 5144 20700
rect 5200 20698 5206 20700
rect 4960 20646 4962 20698
rect 5142 20646 5144 20698
rect 4898 20644 4904 20646
rect 4960 20644 4984 20646
rect 5040 20644 5064 20646
rect 5120 20644 5144 20646
rect 5200 20644 5206 20646
rect 4898 20635 5206 20644
rect 8846 20700 9154 20709
rect 8846 20698 8852 20700
rect 8908 20698 8932 20700
rect 8988 20698 9012 20700
rect 9068 20698 9092 20700
rect 9148 20698 9154 20700
rect 8908 20646 8910 20698
rect 9090 20646 9092 20698
rect 8846 20644 8852 20646
rect 8908 20644 8932 20646
rect 8988 20644 9012 20646
rect 9068 20644 9092 20646
rect 9148 20644 9154 20646
rect 8846 20635 9154 20644
rect 12794 20700 13102 20709
rect 12794 20698 12800 20700
rect 12856 20698 12880 20700
rect 12936 20698 12960 20700
rect 13016 20698 13040 20700
rect 13096 20698 13102 20700
rect 12856 20646 12858 20698
rect 13038 20646 13040 20698
rect 12794 20644 12800 20646
rect 12856 20644 12880 20646
rect 12936 20644 12960 20646
rect 13016 20644 13040 20646
rect 13096 20644 13102 20646
rect 12794 20635 13102 20644
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1688 18970 1716 20402
rect 2924 20156 3232 20165
rect 2924 20154 2930 20156
rect 2986 20154 3010 20156
rect 3066 20154 3090 20156
rect 3146 20154 3170 20156
rect 3226 20154 3232 20156
rect 2986 20102 2988 20154
rect 3168 20102 3170 20154
rect 2924 20100 2930 20102
rect 2986 20100 3010 20102
rect 3066 20100 3090 20102
rect 3146 20100 3170 20102
rect 3226 20100 3232 20102
rect 2924 20091 3232 20100
rect 6872 20156 7180 20165
rect 6872 20154 6878 20156
rect 6934 20154 6958 20156
rect 7014 20154 7038 20156
rect 7094 20154 7118 20156
rect 7174 20154 7180 20156
rect 6934 20102 6936 20154
rect 7116 20102 7118 20154
rect 6872 20100 6878 20102
rect 6934 20100 6958 20102
rect 7014 20100 7038 20102
rect 7094 20100 7118 20102
rect 7174 20100 7180 20102
rect 6872 20091 7180 20100
rect 10820 20156 11128 20165
rect 10820 20154 10826 20156
rect 10882 20154 10906 20156
rect 10962 20154 10986 20156
rect 11042 20154 11066 20156
rect 11122 20154 11128 20156
rect 10882 20102 10884 20154
rect 11064 20102 11066 20154
rect 10820 20100 10826 20102
rect 10882 20100 10906 20102
rect 10962 20100 10986 20102
rect 11042 20100 11066 20102
rect 11122 20100 11128 20102
rect 10820 20091 11128 20100
rect 14768 20156 15076 20165
rect 14768 20154 14774 20156
rect 14830 20154 14854 20156
rect 14910 20154 14934 20156
rect 14990 20154 15014 20156
rect 15070 20154 15076 20156
rect 14830 20102 14832 20154
rect 15012 20102 15014 20154
rect 14768 20100 14774 20102
rect 14830 20100 14854 20102
rect 14910 20100 14934 20102
rect 14990 20100 15014 20102
rect 15070 20100 15076 20102
rect 14768 20091 15076 20100
rect 3330 19952 3386 19961
rect 3330 19887 3386 19896
rect 2924 19068 3232 19077
rect 2924 19066 2930 19068
rect 2986 19066 3010 19068
rect 3066 19066 3090 19068
rect 3146 19066 3170 19068
rect 3226 19066 3232 19068
rect 2986 19014 2988 19066
rect 3168 19014 3170 19066
rect 2924 19012 2930 19014
rect 2986 19012 3010 19014
rect 3066 19012 3090 19014
rect 3146 19012 3170 19014
rect 3226 19012 3232 19014
rect 2924 19003 3232 19012
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2778 18728 2834 18737
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1412 12986 1440 17614
rect 1504 17241 1532 18022
rect 2148 17678 2176 18022
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2332 17338 2360 18702
rect 2778 18663 2834 18672
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1492 17128 1544 17134
rect 1492 17070 1544 17076
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 2320 17128 2372 17134
rect 2320 17070 2372 17076
rect 1400 12980 1452 12986
rect 1400 12922 1452 12928
rect 1504 9722 1532 17070
rect 1964 16726 1992 17070
rect 1952 16720 2004 16726
rect 1952 16662 2004 16668
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1688 14346 1716 16050
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 14958 1808 15438
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1780 14346 1808 14894
rect 1676 14340 1728 14346
rect 1676 14282 1728 14288
rect 1768 14340 1820 14346
rect 1768 14282 1820 14288
rect 1688 13734 1716 14282
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1688 13274 1716 13670
rect 1964 13274 1992 16390
rect 2056 14929 2084 16390
rect 2136 15904 2188 15910
rect 2136 15846 2188 15852
rect 2042 14920 2098 14929
rect 2042 14855 2098 14864
rect 2044 14340 2096 14346
rect 2044 14282 2096 14288
rect 2056 13938 2084 14282
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1688 13258 1808 13274
rect 1964 13258 2084 13274
rect 1688 13252 1820 13258
rect 1688 13246 1768 13252
rect 1964 13252 2096 13258
rect 1964 13246 2044 13252
rect 1768 13194 1820 13200
rect 2044 13194 2096 13200
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1596 11898 1624 12786
rect 2148 12306 2176 15846
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2240 12986 2268 14350
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2332 12782 2360 17070
rect 2424 16454 2452 18226
rect 2792 17882 2820 18663
rect 2924 17980 3232 17989
rect 2924 17978 2930 17980
rect 2986 17978 3010 17980
rect 3066 17978 3090 17980
rect 3146 17978 3170 17980
rect 3226 17978 3232 17980
rect 2986 17926 2988 17978
rect 3168 17926 3170 17978
rect 2924 17924 2930 17926
rect 2986 17924 3010 17926
rect 3066 17924 3090 17926
rect 3146 17924 3170 17926
rect 3226 17924 3232 17926
rect 2924 17915 3232 17924
rect 3344 17882 3372 19887
rect 4898 19612 5206 19621
rect 4898 19610 4904 19612
rect 4960 19610 4984 19612
rect 5040 19610 5064 19612
rect 5120 19610 5144 19612
rect 5200 19610 5206 19612
rect 4960 19558 4962 19610
rect 5142 19558 5144 19610
rect 4898 19556 4904 19558
rect 4960 19556 4984 19558
rect 5040 19556 5064 19558
rect 5120 19556 5144 19558
rect 5200 19556 5206 19558
rect 4898 19547 5206 19556
rect 8846 19612 9154 19621
rect 8846 19610 8852 19612
rect 8908 19610 8932 19612
rect 8988 19610 9012 19612
rect 9068 19610 9092 19612
rect 9148 19610 9154 19612
rect 8908 19558 8910 19610
rect 9090 19558 9092 19610
rect 8846 19556 8852 19558
rect 8908 19556 8932 19558
rect 8988 19556 9012 19558
rect 9068 19556 9092 19558
rect 9148 19556 9154 19558
rect 8846 19547 9154 19556
rect 12794 19612 13102 19621
rect 12794 19610 12800 19612
rect 12856 19610 12880 19612
rect 12936 19610 12960 19612
rect 13016 19610 13040 19612
rect 13096 19610 13102 19612
rect 12856 19558 12858 19610
rect 13038 19558 13040 19610
rect 12794 19556 12800 19558
rect 12856 19556 12880 19558
rect 12936 19556 12960 19558
rect 13016 19556 13040 19558
rect 13096 19556 13102 19558
rect 12794 19547 13102 19556
rect 6872 19068 7180 19077
rect 6872 19066 6878 19068
rect 6934 19066 6958 19068
rect 7014 19066 7038 19068
rect 7094 19066 7118 19068
rect 7174 19066 7180 19068
rect 6934 19014 6936 19066
rect 7116 19014 7118 19066
rect 6872 19012 6878 19014
rect 6934 19012 6958 19014
rect 7014 19012 7038 19014
rect 7094 19012 7118 19014
rect 7174 19012 7180 19014
rect 6872 19003 7180 19012
rect 10820 19068 11128 19077
rect 10820 19066 10826 19068
rect 10882 19066 10906 19068
rect 10962 19066 10986 19068
rect 11042 19066 11066 19068
rect 11122 19066 11128 19068
rect 10882 19014 10884 19066
rect 11064 19014 11066 19066
rect 10820 19012 10826 19014
rect 10882 19012 10906 19014
rect 10962 19012 10986 19014
rect 11042 19012 11066 19014
rect 11122 19012 11128 19014
rect 10820 19003 11128 19012
rect 14768 19068 15076 19077
rect 14768 19066 14774 19068
rect 14830 19066 14854 19068
rect 14910 19066 14934 19068
rect 14990 19066 15014 19068
rect 15070 19066 15076 19068
rect 14830 19014 14832 19066
rect 15012 19014 15014 19066
rect 14768 19012 14774 19014
rect 14830 19012 14854 19014
rect 14910 19012 14934 19014
rect 14990 19012 15014 19014
rect 15070 19012 15076 19014
rect 14768 19003 15076 19012
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 3700 18216 3752 18222
rect 3700 18158 3752 18164
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3332 17604 3384 17610
rect 3332 17546 3384 17552
rect 2924 16892 3232 16901
rect 2924 16890 2930 16892
rect 2986 16890 3010 16892
rect 3066 16890 3090 16892
rect 3146 16890 3170 16892
rect 3226 16890 3232 16892
rect 2986 16838 2988 16890
rect 3168 16838 3170 16890
rect 2924 16836 2930 16838
rect 2986 16836 3010 16838
rect 3066 16836 3090 16838
rect 3146 16836 3170 16838
rect 3226 16836 3232 16838
rect 2924 16827 3232 16836
rect 2504 16516 2556 16522
rect 2504 16458 2556 16464
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2516 12345 2544 16458
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2792 15745 2820 16390
rect 3068 15910 3096 16458
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2924 15804 3232 15813
rect 2924 15802 2930 15804
rect 2986 15802 3010 15804
rect 3066 15802 3090 15804
rect 3146 15802 3170 15804
rect 3226 15802 3232 15804
rect 2986 15750 2988 15802
rect 3168 15750 3170 15802
rect 2924 15748 2930 15750
rect 2986 15748 3010 15750
rect 3066 15748 3090 15750
rect 3146 15748 3170 15750
rect 3226 15748 3232 15750
rect 2778 15736 2834 15745
rect 2924 15739 3232 15748
rect 2778 15671 2834 15680
rect 2924 14716 3232 14725
rect 2924 14714 2930 14716
rect 2986 14714 3010 14716
rect 3066 14714 3090 14716
rect 3146 14714 3170 14716
rect 3226 14714 3232 14716
rect 2986 14662 2988 14714
rect 3168 14662 3170 14714
rect 2924 14660 2930 14662
rect 2986 14660 3010 14662
rect 3066 14660 3090 14662
rect 3146 14660 3170 14662
rect 3226 14660 3232 14662
rect 2924 14651 3232 14660
rect 3344 14249 3372 17546
rect 3712 17338 3740 18158
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3436 15065 3464 15982
rect 3422 15056 3478 15065
rect 3422 14991 3478 15000
rect 3436 14958 3464 14991
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3330 14240 3386 14249
rect 3330 14175 3386 14184
rect 2924 13628 3232 13637
rect 2924 13626 2930 13628
rect 2986 13626 3010 13628
rect 3066 13626 3090 13628
rect 3146 13626 3170 13628
rect 3226 13626 3232 13628
rect 2986 13574 2988 13626
rect 3168 13574 3170 13626
rect 2924 13572 2930 13574
rect 2986 13572 3010 13574
rect 3066 13572 3090 13574
rect 3146 13572 3170 13574
rect 3226 13572 3232 13574
rect 2924 13563 3232 13572
rect 2686 13424 2742 13433
rect 2686 13359 2742 13368
rect 2700 12850 2728 13359
rect 2778 13288 2834 13297
rect 2778 13223 2834 13232
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2792 12442 2820 13223
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 2962 12880 3018 12889
rect 2962 12815 2964 12824
rect 3016 12815 3018 12824
rect 2964 12786 3016 12792
rect 2924 12540 3232 12549
rect 2924 12538 2930 12540
rect 2986 12538 3010 12540
rect 3066 12538 3090 12540
rect 3146 12538 3170 12540
rect 3226 12538 3232 12540
rect 2986 12486 2988 12538
rect 3168 12486 3170 12538
rect 2924 12484 2930 12486
rect 2986 12484 3010 12486
rect 3066 12484 3090 12486
rect 3146 12484 3170 12486
rect 3226 12484 3232 12486
rect 2924 12475 3232 12484
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 3056 12368 3108 12374
rect 2502 12336 2558 12345
rect 2136 12300 2188 12306
rect 3056 12310 3108 12316
rect 2502 12271 2504 12280
rect 2136 12242 2188 12248
rect 2556 12271 2558 12280
rect 2504 12242 2556 12248
rect 2044 12232 2096 12238
rect 2516 12211 2544 12242
rect 2044 12174 2096 12180
rect 2056 12102 2084 12174
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 2056 11676 2084 12038
rect 2136 11688 2188 11694
rect 2056 11648 2136 11676
rect 2136 11630 2188 11636
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2700 11558 2728 11630
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 1676 10600 1728 10606
rect 2516 10577 2544 11018
rect 2792 10713 2820 11630
rect 3068 11626 3096 12310
rect 3344 12306 3372 13126
rect 3528 12753 3556 16934
rect 4344 16720 4396 16726
rect 4344 16662 4396 16668
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3620 15366 3648 15982
rect 3608 15360 3660 15366
rect 3608 15302 3660 15308
rect 3514 12744 3570 12753
rect 3424 12708 3476 12714
rect 3514 12679 3570 12688
rect 3424 12650 3476 12656
rect 3436 12617 3464 12650
rect 3422 12608 3478 12617
rect 3422 12543 3478 12552
rect 3436 12374 3464 12543
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3620 12102 3648 15302
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3804 12850 3832 14214
rect 3896 13569 3924 15982
rect 3988 14006 4016 16390
rect 4356 16046 4384 16662
rect 4540 16250 4568 17614
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4356 15609 4384 15982
rect 4342 15600 4398 15609
rect 4160 15564 4212 15570
rect 4342 15535 4398 15544
rect 4160 15506 4212 15512
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4080 15094 4108 15370
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4080 14006 4108 15030
rect 4172 14618 4200 15506
rect 4356 15502 4384 15535
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4620 15496 4672 15502
rect 4724 15473 4752 16526
rect 4816 15706 4844 18634
rect 4898 18524 5206 18533
rect 4898 18522 4904 18524
rect 4960 18522 4984 18524
rect 5040 18522 5064 18524
rect 5120 18522 5144 18524
rect 5200 18522 5206 18524
rect 4960 18470 4962 18522
rect 5142 18470 5144 18522
rect 4898 18468 4904 18470
rect 4960 18468 4984 18470
rect 5040 18468 5064 18470
rect 5120 18468 5144 18470
rect 5200 18468 5206 18470
rect 4898 18459 5206 18468
rect 8846 18524 9154 18533
rect 8846 18522 8852 18524
rect 8908 18522 8932 18524
rect 8988 18522 9012 18524
rect 9068 18522 9092 18524
rect 9148 18522 9154 18524
rect 8908 18470 8910 18522
rect 9090 18470 9092 18522
rect 8846 18468 8852 18470
rect 8908 18468 8932 18470
rect 8988 18468 9012 18470
rect 9068 18468 9092 18470
rect 9148 18468 9154 18470
rect 8846 18459 9154 18468
rect 12794 18524 13102 18533
rect 12794 18522 12800 18524
rect 12856 18522 12880 18524
rect 12936 18522 12960 18524
rect 13016 18522 13040 18524
rect 13096 18522 13102 18524
rect 12856 18470 12858 18522
rect 13038 18470 13040 18522
rect 12794 18468 12800 18470
rect 12856 18468 12880 18470
rect 12936 18468 12960 18470
rect 13016 18468 13040 18470
rect 13096 18468 13102 18470
rect 12794 18459 13102 18468
rect 6872 17980 7180 17989
rect 6872 17978 6878 17980
rect 6934 17978 6958 17980
rect 7014 17978 7038 17980
rect 7094 17978 7118 17980
rect 7174 17978 7180 17980
rect 6934 17926 6936 17978
rect 7116 17926 7118 17978
rect 6872 17924 6878 17926
rect 6934 17924 6958 17926
rect 7014 17924 7038 17926
rect 7094 17924 7118 17926
rect 7174 17924 7180 17926
rect 6872 17915 7180 17924
rect 10820 17980 11128 17989
rect 10820 17978 10826 17980
rect 10882 17978 10906 17980
rect 10962 17978 10986 17980
rect 11042 17978 11066 17980
rect 11122 17978 11128 17980
rect 10882 17926 10884 17978
rect 11064 17926 11066 17978
rect 10820 17924 10826 17926
rect 10882 17924 10906 17926
rect 10962 17924 10986 17926
rect 11042 17924 11066 17926
rect 11122 17924 11128 17926
rect 10820 17915 11128 17924
rect 14768 17980 15076 17989
rect 14768 17978 14774 17980
rect 14830 17978 14854 17980
rect 14910 17978 14934 17980
rect 14990 17978 15014 17980
rect 15070 17978 15076 17980
rect 14830 17926 14832 17978
rect 15012 17926 15014 17978
rect 14768 17924 14774 17926
rect 14830 17924 14854 17926
rect 14910 17924 14934 17926
rect 14990 17924 15014 17926
rect 15070 17924 15076 17926
rect 14768 17915 15076 17924
rect 4898 17436 5206 17445
rect 4898 17434 4904 17436
rect 4960 17434 4984 17436
rect 5040 17434 5064 17436
rect 5120 17434 5144 17436
rect 5200 17434 5206 17436
rect 4960 17382 4962 17434
rect 5142 17382 5144 17434
rect 4898 17380 4904 17382
rect 4960 17380 4984 17382
rect 5040 17380 5064 17382
rect 5120 17380 5144 17382
rect 5200 17380 5206 17382
rect 4898 17371 5206 17380
rect 8846 17436 9154 17445
rect 8846 17434 8852 17436
rect 8908 17434 8932 17436
rect 8988 17434 9012 17436
rect 9068 17434 9092 17436
rect 9148 17434 9154 17436
rect 8908 17382 8910 17434
rect 9090 17382 9092 17434
rect 8846 17380 8852 17382
rect 8908 17380 8932 17382
rect 8988 17380 9012 17382
rect 9068 17380 9092 17382
rect 9148 17380 9154 17382
rect 8846 17371 9154 17380
rect 12794 17436 13102 17445
rect 12794 17434 12800 17436
rect 12856 17434 12880 17436
rect 12936 17434 12960 17436
rect 13016 17434 13040 17436
rect 13096 17434 13102 17436
rect 12856 17382 12858 17434
rect 13038 17382 13040 17434
rect 12794 17380 12800 17382
rect 12856 17380 12880 17382
rect 12936 17380 12960 17382
rect 13016 17380 13040 17382
rect 13096 17380 13102 17382
rect 12794 17371 13102 17380
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 4898 16348 5206 16357
rect 4898 16346 4904 16348
rect 4960 16346 4984 16348
rect 5040 16346 5064 16348
rect 5120 16346 5144 16348
rect 5200 16346 5206 16348
rect 4960 16294 4962 16346
rect 5142 16294 5144 16346
rect 4898 16292 4904 16294
rect 4960 16292 4984 16294
rect 5040 16292 5064 16294
rect 5120 16292 5144 16294
rect 5200 16292 5206 16294
rect 4898 16283 5206 16292
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5276 15706 5304 15846
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 4620 15438 4672 15444
rect 4710 15464 4766 15473
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 3882 13560 3938 13569
rect 3882 13495 3938 13504
rect 3988 13410 4016 13942
rect 3896 13382 4016 13410
rect 3896 13326 3924 13382
rect 3884 13320 3936 13326
rect 4080 13274 4108 13942
rect 3884 13262 3936 13268
rect 3988 13246 4108 13274
rect 4264 13258 4292 14962
rect 4252 13252 4304 13258
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3988 12442 4016 13246
rect 4252 13194 4304 13200
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 2924 11452 3232 11461
rect 2924 11450 2930 11452
rect 2986 11450 3010 11452
rect 3066 11450 3090 11452
rect 3146 11450 3170 11452
rect 3226 11450 3232 11452
rect 2986 11398 2988 11450
rect 3168 11398 3170 11450
rect 2924 11396 2930 11398
rect 2986 11396 3010 11398
rect 3066 11396 3090 11398
rect 3146 11396 3170 11398
rect 3226 11396 3232 11398
rect 2924 11387 3232 11396
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 2778 10704 2834 10713
rect 2778 10639 2834 10648
rect 1676 10542 1728 10548
rect 2502 10568 2558 10577
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1492 9716 1544 9722
rect 1492 9658 1544 9664
rect 1306 9480 1362 9489
rect 1306 9415 1362 9424
rect 1320 3369 1348 9415
rect 1504 9081 1532 9658
rect 1490 9072 1546 9081
rect 1596 9042 1624 9862
rect 1688 9178 1716 10542
rect 2502 10503 2558 10512
rect 2924 10364 3232 10373
rect 2924 10362 2930 10364
rect 2986 10362 3010 10364
rect 3066 10362 3090 10364
rect 3146 10362 3170 10364
rect 3226 10362 3232 10364
rect 2986 10310 2988 10362
rect 3168 10310 3170 10362
rect 2924 10308 2930 10310
rect 2986 10308 3010 10310
rect 3066 10308 3090 10310
rect 3146 10308 3170 10310
rect 3226 10308 3232 10310
rect 2924 10299 3232 10308
rect 3436 10169 3464 11086
rect 3528 10810 3556 11630
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3422 10160 3478 10169
rect 3422 10095 3478 10104
rect 1766 10024 1822 10033
rect 1766 9959 1768 9968
rect 1820 9959 1822 9968
rect 3332 9988 3384 9994
rect 1768 9930 1820 9936
rect 3332 9930 3384 9936
rect 2924 9276 3232 9285
rect 2924 9274 2930 9276
rect 2986 9274 3010 9276
rect 3066 9274 3090 9276
rect 3146 9274 3170 9276
rect 3226 9274 3232 9276
rect 2986 9222 2988 9274
rect 3168 9222 3170 9274
rect 2924 9220 2930 9222
rect 2986 9220 3010 9222
rect 3066 9220 3090 9222
rect 3146 9220 3170 9222
rect 3226 9220 3232 9222
rect 2924 9211 3232 9220
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 1490 9007 1546 9016
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 6866 1440 8366
rect 1596 7750 1624 8978
rect 1688 8838 1716 9114
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 2042 7848 2098 7857
rect 1676 7812 1728 7818
rect 2042 7783 2098 7792
rect 1676 7754 1728 7760
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 7002 1532 7346
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1398 6760 1454 6769
rect 1398 6695 1454 6704
rect 1412 4690 1440 6695
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1504 4593 1532 6258
rect 1596 6225 1624 7686
rect 1582 6216 1638 6225
rect 1582 6151 1638 6160
rect 1490 4584 1546 4593
rect 1490 4519 1546 4528
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 1412 3777 1440 4014
rect 1398 3768 1454 3777
rect 1398 3703 1454 3712
rect 1306 3360 1362 3369
rect 1306 3295 1362 3304
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 2281 1440 2382
rect 1398 2272 1454 2281
rect 1398 2207 1454 2216
rect 1400 1352 1452 1358
rect 1400 1294 1452 1300
rect 1412 785 1440 1294
rect 1504 1222 1532 4519
rect 1596 3058 1624 6151
rect 1688 4690 1716 7754
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1858 7304 1914 7313
rect 1780 5778 1808 7278
rect 1858 7239 1914 7248
rect 1872 6390 1900 7239
rect 1860 6384 1912 6390
rect 1860 6326 1912 6332
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1780 4146 1808 5714
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1674 4040 1730 4049
rect 1674 3975 1730 3984
rect 1688 3534 1716 3975
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1872 3126 1900 6326
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1964 2650 1992 6258
rect 2056 3602 2084 7783
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2148 3398 2176 7142
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2240 3534 2268 4422
rect 2332 3738 2360 8842
rect 2976 8838 3004 9114
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2686 8528 2742 8537
rect 2686 8463 2742 8472
rect 2700 7750 2728 8463
rect 2924 8188 3232 8197
rect 2924 8186 2930 8188
rect 2986 8186 3010 8188
rect 3066 8186 3090 8188
rect 3146 8186 3170 8188
rect 3226 8186 3232 8188
rect 2986 8134 2988 8186
rect 3168 8134 3170 8186
rect 2924 8132 2930 8134
rect 2986 8132 3010 8134
rect 3066 8132 3090 8134
rect 3146 8132 3170 8134
rect 3226 8132 3232 8134
rect 2924 8123 3232 8132
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2424 6390 2452 7278
rect 2792 6916 2820 7822
rect 3252 7478 3280 7890
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3068 7206 3096 7346
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 2924 7100 3232 7109
rect 2924 7098 2930 7100
rect 2986 7098 3010 7100
rect 3066 7098 3090 7100
rect 3146 7098 3170 7100
rect 3226 7098 3232 7100
rect 2986 7046 2988 7098
rect 3168 7046 3170 7098
rect 2924 7044 2930 7046
rect 2986 7044 3010 7046
rect 3066 7044 3090 7046
rect 3146 7044 3170 7046
rect 3226 7044 3232 7046
rect 2924 7035 3232 7044
rect 2872 6928 2924 6934
rect 2792 6888 2872 6916
rect 2872 6870 2924 6876
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2412 6384 2464 6390
rect 2792 6361 2820 6394
rect 2412 6326 2464 6332
rect 2778 6352 2834 6361
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2424 3194 2452 6326
rect 3160 6322 3188 6802
rect 2778 6287 2834 6296
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2924 6012 3232 6021
rect 2924 6010 2930 6012
rect 2986 6010 3010 6012
rect 3066 6010 3090 6012
rect 3146 6010 3170 6012
rect 3226 6010 3232 6012
rect 2986 5958 2988 6010
rect 3168 5958 3170 6010
rect 2924 5956 2930 5958
rect 2986 5956 3010 5958
rect 3066 5956 3090 5958
rect 3146 5956 3170 5958
rect 3226 5956 3232 5958
rect 2924 5947 3232 5956
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2608 5574 2636 5646
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2516 4078 2544 5170
rect 2608 5166 2636 5510
rect 3054 5400 3110 5409
rect 3054 5335 3110 5344
rect 3068 5234 3096 5335
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2226 3088 2282 3097
rect 2516 3058 2544 4014
rect 2226 3023 2228 3032
rect 2280 3023 2282 3032
rect 2504 3052 2556 3058
rect 2228 2994 2280 3000
rect 2504 2994 2556 3000
rect 2608 2774 2636 5102
rect 3068 5012 3096 5170
rect 3252 5137 3280 5170
rect 3238 5128 3294 5137
rect 3238 5063 3294 5072
rect 2859 4984 3096 5012
rect 2859 4808 2887 4984
rect 2924 4924 3232 4933
rect 2924 4922 2930 4924
rect 2986 4922 3010 4924
rect 3066 4922 3090 4924
rect 3146 4922 3170 4924
rect 3226 4922 3232 4924
rect 2986 4870 2988 4922
rect 3168 4870 3170 4922
rect 2924 4868 2930 4870
rect 2986 4868 3010 4870
rect 3066 4868 3090 4870
rect 3146 4868 3170 4870
rect 3226 4868 3232 4870
rect 2924 4859 3232 4868
rect 3056 4820 3108 4826
rect 2859 4780 2912 4808
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2700 3670 2728 4558
rect 2884 4282 2912 4780
rect 3056 4762 3108 4768
rect 3068 4729 3096 4762
rect 3054 4720 3110 4729
rect 3054 4655 3110 4664
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2870 4176 2926 4185
rect 2870 4111 2872 4120
rect 2924 4111 2926 4120
rect 2872 4082 2924 4088
rect 2884 3924 2912 4082
rect 2976 4078 3004 4218
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2859 3896 2912 3924
rect 2859 3720 2887 3896
rect 2924 3836 3232 3845
rect 2924 3834 2930 3836
rect 2986 3834 3010 3836
rect 3066 3834 3090 3836
rect 3146 3834 3170 3836
rect 3226 3834 3232 3836
rect 2986 3782 2988 3834
rect 3168 3782 3170 3834
rect 2924 3780 2930 3782
rect 2986 3780 3010 3782
rect 3066 3780 3090 3782
rect 3146 3780 3170 3782
rect 3226 3780 3232 3782
rect 2924 3771 3232 3780
rect 2859 3692 2912 3720
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2778 3632 2834 3641
rect 2884 3618 2912 3692
rect 2884 3590 3096 3618
rect 2778 3567 2834 3576
rect 2608 2746 2728 2774
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2700 2582 2728 2746
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2056 1970 2084 2450
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2700 1970 2728 2382
rect 2044 1964 2096 1970
rect 2044 1906 2096 1912
rect 2688 1964 2740 1970
rect 2688 1906 2740 1912
rect 2792 1902 2820 3567
rect 3068 3534 3096 3590
rect 2964 3528 3016 3534
rect 2962 3496 2964 3505
rect 3056 3528 3108 3534
rect 3016 3496 3018 3505
rect 3056 3470 3108 3476
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 2962 3431 3018 3440
rect 3160 3369 3188 3470
rect 3146 3360 3202 3369
rect 3146 3295 3202 3304
rect 3344 3194 3372 9930
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 8906 3464 9318
rect 3528 8974 3556 10474
rect 3712 10266 3740 11630
rect 3804 11354 3832 12174
rect 4172 11898 4200 12718
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4264 11665 4292 13194
rect 4250 11656 4306 11665
rect 4250 11591 4306 11600
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 4264 10742 4292 11591
rect 4356 11150 4384 15438
rect 4632 14906 4660 15438
rect 4710 15399 4766 15408
rect 4898 15260 5206 15269
rect 4898 15258 4904 15260
rect 4960 15258 4984 15260
rect 5040 15258 5064 15260
rect 5120 15258 5144 15260
rect 5200 15258 5206 15260
rect 4960 15206 4962 15258
rect 5142 15206 5144 15258
rect 4898 15204 4904 15206
rect 4960 15204 4984 15206
rect 5040 15204 5064 15206
rect 5120 15204 5144 15206
rect 5200 15204 5206 15206
rect 4898 15195 5206 15204
rect 5356 14952 5408 14958
rect 4632 14878 4752 14906
rect 5356 14894 5408 14900
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4540 14618 4568 14758
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 4448 12850 4476 14282
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 4448 11830 4476 12786
rect 4632 12306 4660 14758
rect 4724 12889 4752 14878
rect 4898 14172 5206 14181
rect 4898 14170 4904 14172
rect 4960 14170 4984 14172
rect 5040 14170 5064 14172
rect 5120 14170 5144 14172
rect 5200 14170 5206 14172
rect 4960 14118 4962 14170
rect 5142 14118 5144 14170
rect 4898 14116 4904 14118
rect 4960 14116 4984 14118
rect 5040 14116 5064 14118
rect 5120 14116 5144 14118
rect 5200 14116 5206 14118
rect 4898 14107 5206 14116
rect 5368 13274 5396 14894
rect 5460 14550 5488 16050
rect 5722 15600 5778 15609
rect 5722 15535 5724 15544
rect 5776 15535 5778 15544
rect 5724 15506 5776 15512
rect 5828 15473 5856 16050
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 5814 15464 5870 15473
rect 5814 15399 5870 15408
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5446 14104 5502 14113
rect 5446 14039 5502 14048
rect 5460 13870 5488 14039
rect 5552 13938 5580 14758
rect 5736 13977 5764 14962
rect 5828 14278 5856 15302
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 6012 14385 6040 14962
rect 5998 14376 6054 14385
rect 5998 14311 6054 14320
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 5722 13968 5778 13977
rect 5540 13932 5592 13938
rect 5592 13892 5672 13920
rect 5722 13903 5778 13912
rect 5908 13932 5960 13938
rect 5540 13874 5592 13880
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5460 13394 5488 13670
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5368 13246 5580 13274
rect 4898 13084 5206 13093
rect 4898 13082 4904 13084
rect 4960 13082 4984 13084
rect 5040 13082 5064 13084
rect 5120 13082 5144 13084
rect 5200 13082 5206 13084
rect 4960 13030 4962 13082
rect 5142 13030 5144 13082
rect 4898 13028 4904 13030
rect 4960 13028 4984 13030
rect 5040 13028 5064 13030
rect 5120 13028 5144 13030
rect 5200 13028 5206 13030
rect 4898 13019 5206 13028
rect 4710 12880 4766 12889
rect 4710 12815 4766 12824
rect 5552 12753 5580 13246
rect 5644 12866 5672 13892
rect 5908 13874 5960 13880
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5736 12986 5764 13806
rect 5920 13802 5948 13874
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5644 12838 5764 12866
rect 5538 12744 5594 12753
rect 5538 12679 5594 12688
rect 4986 12608 5042 12617
rect 4986 12543 5042 12552
rect 5000 12306 5028 12543
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4724 11014 4752 12174
rect 4898 11996 5206 12005
rect 4898 11994 4904 11996
rect 4960 11994 4984 11996
rect 5040 11994 5064 11996
rect 5120 11994 5144 11996
rect 5200 11994 5206 11996
rect 4960 11942 4962 11994
rect 5142 11942 5144 11994
rect 4898 11940 4904 11942
rect 4960 11940 4984 11942
rect 5040 11940 5064 11942
rect 5120 11940 5144 11942
rect 5200 11940 5206 11942
rect 4898 11931 5206 11940
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5460 11218 5488 11698
rect 5552 11626 5580 12679
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5644 11354 5672 12174
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4898 10908 5206 10917
rect 4898 10906 4904 10908
rect 4960 10906 4984 10908
rect 5040 10906 5064 10908
rect 5120 10906 5144 10908
rect 5200 10906 5206 10908
rect 4960 10854 4962 10906
rect 5142 10854 5144 10906
rect 4898 10852 4904 10854
rect 4960 10852 4984 10854
rect 5040 10852 5064 10854
rect 5120 10852 5144 10854
rect 5200 10852 5206 10854
rect 4898 10843 5206 10852
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 4080 10033 4108 10678
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3516 8968 3568 8974
rect 3514 8936 3516 8945
rect 3568 8936 3570 8945
rect 3424 8900 3476 8906
rect 3514 8871 3570 8880
rect 3424 8842 3476 8848
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3528 8401 3556 8434
rect 3514 8392 3570 8401
rect 3514 8327 3570 8336
rect 3422 7984 3478 7993
rect 3422 7919 3478 7928
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 3160 2922 3188 3062
rect 3148 2916 3200 2922
rect 3148 2858 3200 2864
rect 2924 2748 3232 2757
rect 2924 2746 2930 2748
rect 2986 2746 3010 2748
rect 3066 2746 3090 2748
rect 3146 2746 3170 2748
rect 3226 2746 3232 2748
rect 2986 2694 2988 2746
rect 3168 2694 3170 2746
rect 2924 2692 2930 2694
rect 2986 2692 3010 2694
rect 3066 2692 3090 2694
rect 3146 2692 3170 2694
rect 3226 2692 3232 2694
rect 2924 2683 3232 2692
rect 3436 2038 3464 7919
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7546 3556 7686
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3528 7206 3556 7346
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 6254 3556 7142
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3528 5302 3556 6054
rect 3620 5370 3648 9862
rect 4264 9722 4292 10406
rect 4908 10062 4936 10678
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3516 5296 3568 5302
rect 3516 5238 3568 5244
rect 3606 4312 3662 4321
rect 3606 4247 3662 4256
rect 3620 4214 3648 4247
rect 3608 4208 3660 4214
rect 3608 4150 3660 4156
rect 3620 2106 3648 4150
rect 3712 3670 3740 9454
rect 3804 8294 3832 9454
rect 3804 8266 3924 8294
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3804 6662 3832 7822
rect 3896 7478 3924 8266
rect 3988 8265 4016 9590
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 3974 8256 4030 8265
rect 3974 8191 4030 8200
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3804 5846 3832 6122
rect 3896 6089 3924 6870
rect 3882 6080 3938 6089
rect 3882 6015 3938 6024
rect 3792 5840 3844 5846
rect 3988 5817 4016 7346
rect 4080 7002 4108 7754
rect 4172 7041 4200 9522
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 4264 9178 4292 9386
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4264 7449 4292 8026
rect 4250 7440 4306 7449
rect 4250 7375 4306 7384
rect 4158 7032 4214 7041
rect 4068 6996 4120 7002
rect 4158 6967 4214 6976
rect 4068 6938 4120 6944
rect 4160 6928 4212 6934
rect 4066 6896 4122 6905
rect 4160 6870 4212 6876
rect 4066 6831 4068 6840
rect 4120 6831 4122 6840
rect 4068 6802 4120 6808
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3792 5782 3844 5788
rect 3974 5808 4030 5817
rect 3974 5743 4030 5752
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3804 5273 3832 5646
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 3988 5352 4016 5578
rect 3896 5324 4016 5352
rect 3790 5264 3846 5273
rect 3790 5199 3846 5208
rect 3896 4010 3924 5324
rect 3974 5264 4030 5273
rect 3974 5199 3976 5208
rect 4028 5199 4030 5208
rect 3976 5170 4028 5176
rect 4080 5098 4108 6598
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 4066 4856 4122 4865
rect 4066 4791 4068 4800
rect 4120 4791 4122 4800
rect 4068 4762 4120 4768
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 3976 4072 4028 4078
rect 3974 4040 3976 4049
rect 4028 4040 4030 4049
rect 3884 4004 3936 4010
rect 3974 3975 4030 3984
rect 3884 3946 3936 3952
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3896 3534 3924 3946
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 4080 3398 4108 4558
rect 4172 4486 4200 6870
rect 4264 6798 4292 7375
rect 4448 6866 4476 9930
rect 4898 9820 5206 9829
rect 4898 9818 4904 9820
rect 4960 9818 4984 9820
rect 5040 9818 5064 9820
rect 5120 9818 5144 9820
rect 5200 9818 5206 9820
rect 4960 9766 4962 9818
rect 5142 9766 5144 9818
rect 4898 9764 4904 9766
rect 4960 9764 4984 9766
rect 5040 9764 5064 9766
rect 5120 9764 5144 9766
rect 5200 9764 5206 9766
rect 4898 9755 5206 9764
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4448 6390 4476 6598
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4264 5642 4292 6258
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4264 5234 4292 5578
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4264 4214 4292 5170
rect 4356 4554 4384 6190
rect 4448 4690 4476 6326
rect 4540 5914 4568 8978
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4540 5166 4568 5714
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4540 4214 4568 4762
rect 4632 4622 4660 8978
rect 4710 8528 4766 8537
rect 4710 8463 4766 8472
rect 4724 8430 4752 8463
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 8090 4752 8230
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4710 7984 4766 7993
rect 4710 7919 4766 7928
rect 4724 7274 4752 7919
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4710 6760 4766 6769
rect 4710 6695 4766 6704
rect 4724 6390 4752 6695
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4816 5030 4844 9318
rect 4898 8732 5206 8741
rect 4898 8730 4904 8732
rect 4960 8730 4984 8732
rect 5040 8730 5064 8732
rect 5120 8730 5144 8732
rect 5200 8730 5206 8732
rect 4960 8678 4962 8730
rect 5142 8678 5144 8730
rect 4898 8676 4904 8678
rect 4960 8676 4984 8678
rect 5040 8676 5064 8678
rect 5120 8676 5144 8678
rect 5200 8676 5206 8678
rect 4898 8667 5206 8676
rect 5264 8560 5316 8566
rect 5078 8528 5134 8537
rect 5264 8502 5316 8508
rect 5078 8463 5134 8472
rect 5092 8362 5120 8463
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 5092 7750 5120 8298
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4898 7644 5206 7653
rect 4898 7642 4904 7644
rect 4960 7642 4984 7644
rect 5040 7642 5064 7644
rect 5120 7642 5144 7644
rect 5200 7642 5206 7644
rect 4960 7590 4962 7642
rect 5142 7590 5144 7642
rect 4898 7588 4904 7590
rect 4960 7588 4984 7590
rect 5040 7588 5064 7590
rect 5120 7588 5144 7590
rect 5200 7588 5206 7590
rect 4898 7579 5206 7588
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 6662 5028 7142
rect 5170 7032 5226 7041
rect 5170 6967 5172 6976
rect 5224 6967 5226 6976
rect 5172 6938 5224 6944
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4898 6556 5206 6565
rect 4898 6554 4904 6556
rect 4960 6554 4984 6556
rect 5040 6554 5064 6556
rect 5120 6554 5144 6556
rect 5200 6554 5206 6556
rect 4960 6502 4962 6554
rect 5142 6502 5144 6554
rect 4898 6500 4904 6502
rect 4960 6500 4984 6502
rect 5040 6500 5064 6502
rect 5120 6500 5144 6502
rect 5200 6500 5206 6502
rect 4898 6491 5206 6500
rect 4988 6452 5040 6458
rect 5040 6412 5120 6440
rect 4988 6394 5040 6400
rect 5092 6322 5120 6412
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5000 5817 5028 6190
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 4986 5808 5042 5817
rect 4986 5743 5042 5752
rect 5092 5681 5120 6122
rect 5078 5672 5134 5681
rect 5078 5607 5134 5616
rect 4898 5468 5206 5477
rect 4898 5466 4904 5468
rect 4960 5466 4984 5468
rect 5040 5466 5064 5468
rect 5120 5466 5144 5468
rect 5200 5466 5206 5468
rect 4960 5414 4962 5466
rect 5142 5414 5144 5466
rect 4898 5412 4904 5414
rect 4960 5412 4984 5414
rect 5040 5412 5064 5414
rect 5120 5412 5144 5414
rect 5200 5412 5206 5414
rect 4898 5403 5206 5412
rect 4712 5024 4764 5030
rect 4710 4992 4712 5001
rect 4804 5024 4856 5030
rect 4764 4992 4766 5001
rect 4804 4966 4856 4972
rect 4710 4927 4766 4936
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4632 4146 4660 4558
rect 5000 4554 5028 4626
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 4898 4380 5206 4389
rect 4898 4378 4904 4380
rect 4960 4378 4984 4380
rect 5040 4378 5064 4380
rect 5120 4378 5144 4380
rect 5200 4378 5206 4380
rect 4960 4326 4962 4378
rect 5142 4326 5144 4378
rect 4898 4324 4904 4326
rect 4960 4324 4984 4326
rect 5040 4324 5064 4326
rect 5120 4324 5144 4326
rect 5200 4324 5206 4326
rect 4898 4315 5206 4324
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4356 3738 4384 3878
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 5092 3602 5120 4082
rect 5276 4010 5304 8502
rect 5368 6458 5396 10610
rect 5460 10606 5488 11154
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5552 10130 5580 11086
rect 5630 10704 5686 10713
rect 5630 10639 5686 10648
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5460 8294 5488 8842
rect 5460 8266 5580 8294
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5368 5710 5396 6258
rect 5356 5704 5408 5710
rect 5460 5681 5488 7754
rect 5552 7721 5580 8266
rect 5644 7886 5672 10639
rect 5736 8129 5764 12838
rect 5920 11898 5948 13738
rect 6012 13530 6040 14214
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6104 13376 6132 15846
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6196 14618 6224 15438
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6288 13802 6316 17002
rect 6872 16892 7180 16901
rect 6872 16890 6878 16892
rect 6934 16890 6958 16892
rect 7014 16890 7038 16892
rect 7094 16890 7118 16892
rect 7174 16890 7180 16892
rect 6934 16838 6936 16890
rect 7116 16838 7118 16890
rect 6872 16836 6878 16838
rect 6934 16836 6958 16838
rect 7014 16836 7038 16838
rect 7094 16836 7118 16838
rect 7174 16836 7180 16838
rect 6872 16827 7180 16836
rect 10820 16892 11128 16901
rect 10820 16890 10826 16892
rect 10882 16890 10906 16892
rect 10962 16890 10986 16892
rect 11042 16890 11066 16892
rect 11122 16890 11128 16892
rect 10882 16838 10884 16890
rect 11064 16838 11066 16890
rect 10820 16836 10826 16838
rect 10882 16836 10906 16838
rect 10962 16836 10986 16838
rect 11042 16836 11066 16838
rect 11122 16836 11128 16838
rect 10820 16827 11128 16836
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6366 14920 6422 14929
rect 6366 14855 6368 14864
rect 6420 14855 6422 14864
rect 6368 14826 6420 14832
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 6104 13348 6224 13376
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5722 8120 5778 8129
rect 5722 8055 5778 8064
rect 5828 8004 5856 11562
rect 5920 10742 5948 11834
rect 6104 11082 6132 13194
rect 6196 12238 6224 13348
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6196 11762 6224 12174
rect 6380 12170 6408 14214
rect 6472 13326 6500 15574
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6564 13258 6592 14486
rect 6748 14090 6776 16458
rect 8846 16348 9154 16357
rect 8846 16346 8852 16348
rect 8908 16346 8932 16348
rect 8988 16346 9012 16348
rect 9068 16346 9092 16348
rect 9148 16346 9154 16348
rect 8908 16294 8910 16346
rect 9090 16294 9092 16346
rect 8846 16292 8852 16294
rect 8908 16292 8932 16294
rect 8988 16292 9012 16294
rect 9068 16292 9092 16294
rect 9148 16292 9154 16294
rect 8846 16283 9154 16292
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 6872 15804 7180 15813
rect 6872 15802 6878 15804
rect 6934 15802 6958 15804
rect 7014 15802 7038 15804
rect 7094 15802 7118 15804
rect 7174 15802 7180 15804
rect 6934 15750 6936 15802
rect 7116 15750 7118 15802
rect 6872 15748 6878 15750
rect 6934 15748 6958 15750
rect 7014 15748 7038 15750
rect 7094 15748 7118 15750
rect 7174 15748 7180 15750
rect 6872 15739 7180 15748
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7024 14890 7052 14962
rect 7116 14929 7144 14962
rect 7102 14920 7158 14929
rect 7012 14884 7064 14890
rect 7102 14855 7158 14864
rect 7012 14826 7064 14832
rect 6872 14716 7180 14725
rect 6872 14714 6878 14716
rect 6934 14714 6958 14716
rect 7014 14714 7038 14716
rect 7094 14714 7118 14716
rect 7174 14714 7180 14716
rect 6934 14662 6936 14714
rect 7116 14662 7118 14714
rect 6872 14660 6878 14662
rect 6934 14660 6958 14662
rect 7014 14660 7038 14662
rect 7094 14660 7118 14662
rect 7174 14660 7180 14662
rect 6872 14651 7180 14660
rect 7208 14482 7236 15370
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 6748 14074 6868 14090
rect 6748 14068 6880 14074
rect 6748 14062 6828 14068
rect 6828 14010 6880 14016
rect 6932 13870 6960 14418
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6748 13433 6776 13738
rect 7208 13734 7236 14282
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 6872 13628 7180 13637
rect 6872 13626 6878 13628
rect 6934 13626 6958 13628
rect 7014 13626 7038 13628
rect 7094 13626 7118 13628
rect 7174 13626 7180 13628
rect 6934 13574 6936 13626
rect 7116 13574 7118 13626
rect 6872 13572 6878 13574
rect 6934 13572 6958 13574
rect 7014 13572 7038 13574
rect 7094 13572 7118 13574
rect 7174 13572 7180 13574
rect 6872 13563 7180 13572
rect 6734 13424 6790 13433
rect 6734 13359 6790 13368
rect 6552 13252 6604 13258
rect 6748 13240 6776 13359
rect 7208 13326 7236 13670
rect 7300 13530 7328 14350
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 6920 13252 6972 13258
rect 6748 13212 6920 13240
rect 6552 13194 6604 13200
rect 6920 13194 6972 13200
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 6472 12050 6500 12106
rect 6288 12022 6500 12050
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 6288 10538 6316 12022
rect 6564 10810 6592 12922
rect 6872 12540 7180 12549
rect 6872 12538 6878 12540
rect 6934 12538 6958 12540
rect 7014 12538 7038 12540
rect 7094 12538 7118 12540
rect 7174 12538 7180 12540
rect 6934 12486 6936 12538
rect 7116 12486 7118 12538
rect 6872 12484 6878 12486
rect 6934 12484 6958 12486
rect 7014 12484 7038 12486
rect 7094 12484 7118 12486
rect 7174 12484 7180 12486
rect 6872 12475 7180 12484
rect 6734 12336 6790 12345
rect 6734 12271 6790 12280
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6656 11529 6684 11766
rect 6642 11520 6698 11529
rect 6642 11455 6698 11464
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6368 10736 6420 10742
rect 6368 10678 6420 10684
rect 6380 10606 6408 10678
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 6380 10266 6408 10542
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5920 8838 5948 9658
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6104 8974 6132 9454
rect 6092 8968 6144 8974
rect 6090 8936 6092 8945
rect 6144 8936 6146 8945
rect 6090 8871 6146 8880
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5736 7976 5856 8004
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5736 7732 5764 7976
rect 5920 7750 5948 8774
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 6012 7954 6040 8298
rect 6196 8129 6224 9998
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6288 9042 6316 9930
rect 6380 9518 6408 10202
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6182 8120 6238 8129
rect 6182 8055 6238 8064
rect 6288 8004 6316 8842
rect 6380 8129 6408 9454
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6564 9178 6592 9318
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6366 8120 6422 8129
rect 6366 8055 6422 8064
rect 6104 7976 6316 8004
rect 6366 7984 6422 7993
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5908 7744 5960 7750
rect 5538 7712 5594 7721
rect 5538 7647 5594 7656
rect 5676 7704 5764 7732
rect 5828 7704 5908 7732
rect 5676 7562 5704 7704
rect 5644 7534 5704 7562
rect 5644 7410 5672 7534
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5828 7290 5856 7704
rect 5908 7686 5960 7692
rect 5906 7576 5962 7585
rect 6104 7562 6132 7976
rect 6366 7919 6422 7928
rect 6380 7886 6408 7919
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6288 7732 6316 7822
rect 6368 7744 6420 7750
rect 6288 7704 6368 7732
rect 6368 7686 6420 7692
rect 6104 7534 6224 7562
rect 5906 7511 5962 7520
rect 5920 7410 5948 7511
rect 5908 7404 5960 7410
rect 6196 7398 6224 7534
rect 6472 7460 6500 9114
rect 6550 9072 6606 9081
rect 6550 9007 6606 9016
rect 6564 8430 6592 9007
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6380 7432 6500 7460
rect 6380 7398 6408 7432
rect 5908 7346 5960 7352
rect 6104 7370 6224 7398
rect 6288 7370 6408 7398
rect 5630 7168 5686 7177
rect 5630 7103 5686 7112
rect 5644 7002 5672 7103
rect 5736 7018 5764 7278
rect 5828 7262 5948 7290
rect 5632 6996 5684 7002
rect 5736 6990 5859 7018
rect 5632 6938 5684 6944
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5630 6896 5686 6905
rect 5552 6610 5580 6870
rect 5831 6882 5859 6990
rect 5686 6854 5764 6882
rect 5630 6831 5686 6840
rect 5552 6582 5672 6610
rect 5644 6322 5672 6582
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5356 5646 5408 5652
rect 5446 5672 5502 5681
rect 5446 5607 5502 5616
rect 5644 5409 5672 5714
rect 5354 5400 5410 5409
rect 5630 5400 5686 5409
rect 5354 5335 5356 5344
rect 5408 5335 5410 5344
rect 5540 5364 5592 5370
rect 5356 5306 5408 5312
rect 5630 5335 5686 5344
rect 5540 5306 5592 5312
rect 5552 5234 5580 5306
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4486 5396 4966
rect 5552 4758 5580 5170
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5644 3913 5672 5335
rect 5736 5234 5764 6854
rect 5828 6854 5859 6882
rect 5828 6730 5856 6854
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5814 6624 5870 6633
rect 5814 6559 5870 6568
rect 5828 6458 5856 6559
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5814 5536 5870 5545
rect 5814 5471 5870 5480
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5828 4826 5856 5471
rect 5920 5166 5948 7262
rect 6104 7002 6132 7370
rect 6288 7324 6316 7370
rect 6196 7296 6316 7324
rect 6460 7336 6512 7342
rect 6000 6996 6052 7002
rect 6092 6996 6144 7002
rect 6052 6956 6092 6984
rect 6000 6938 6052 6944
rect 6092 6938 6144 6944
rect 6196 6848 6224 7296
rect 6564 7324 6592 8230
rect 6656 7392 6684 9318
rect 6748 8498 6776 12271
rect 6826 12200 6882 12209
rect 6826 12135 6882 12144
rect 6840 12102 6868 12135
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6872 11452 7180 11461
rect 6872 11450 6878 11452
rect 6934 11450 6958 11452
rect 7014 11450 7038 11452
rect 7094 11450 7118 11452
rect 7174 11450 7180 11452
rect 6934 11398 6936 11450
rect 7116 11398 7118 11450
rect 6872 11396 6878 11398
rect 6934 11396 6958 11398
rect 7014 11396 7038 11398
rect 7094 11396 7118 11398
rect 7174 11396 7180 11398
rect 6872 11387 7180 11396
rect 7208 11150 7236 13262
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 6872 10364 7180 10373
rect 6872 10362 6878 10364
rect 6934 10362 6958 10364
rect 7014 10362 7038 10364
rect 7094 10362 7118 10364
rect 7174 10362 7180 10364
rect 6934 10310 6936 10362
rect 7116 10310 7118 10362
rect 6872 10308 6878 10310
rect 6934 10308 6958 10310
rect 7014 10308 7038 10310
rect 7094 10308 7118 10310
rect 7174 10308 7180 10310
rect 6872 10299 7180 10308
rect 7300 10266 7328 13194
rect 7392 11354 7420 15438
rect 7654 15056 7710 15065
rect 7654 14991 7710 15000
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13138 7512 14214
rect 7562 14104 7618 14113
rect 7562 14039 7618 14048
rect 7576 13326 7604 14039
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7484 13110 7604 13138
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7484 11665 7512 11698
rect 7470 11656 7526 11665
rect 7470 11591 7526 11600
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7484 11150 7512 11494
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7484 10538 7512 10950
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6872 9276 7180 9285
rect 6872 9274 6878 9276
rect 6934 9274 6958 9276
rect 7014 9274 7038 9276
rect 7094 9274 7118 9276
rect 7174 9274 7180 9276
rect 6934 9222 6936 9274
rect 7116 9222 7118 9274
rect 6872 9220 6878 9222
rect 6934 9220 6958 9222
rect 7014 9220 7038 9222
rect 7094 9220 7118 9222
rect 7174 9220 7180 9222
rect 6872 9211 7180 9220
rect 7102 8936 7158 8945
rect 7102 8871 7158 8880
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6840 8537 6868 8570
rect 6826 8528 6882 8537
rect 6736 8492 6788 8498
rect 7116 8498 7144 8871
rect 6826 8463 6882 8472
rect 7104 8492 7156 8498
rect 6736 8434 6788 8440
rect 7104 8434 7156 8440
rect 6872 8188 7180 8197
rect 6872 8186 6878 8188
rect 6934 8186 6958 8188
rect 7014 8186 7038 8188
rect 7094 8186 7118 8188
rect 7174 8186 7180 8188
rect 6934 8134 6936 8186
rect 7116 8134 7118 8186
rect 6872 8132 6878 8134
rect 6934 8132 6958 8134
rect 7014 8132 7038 8134
rect 7094 8132 7118 8134
rect 7174 8132 7180 8134
rect 6872 8123 7180 8132
rect 7104 8016 7156 8022
rect 7102 7984 7104 7993
rect 7156 7984 7158 7993
rect 6828 7948 6880 7954
rect 7102 7919 7158 7928
rect 6828 7890 6880 7896
rect 6840 7449 6868 7890
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 7478 7052 7686
rect 7116 7585 7144 7822
rect 7102 7576 7158 7585
rect 7208 7546 7236 9522
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7300 7750 7328 9046
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7102 7511 7158 7520
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7012 7472 7064 7478
rect 6826 7440 6882 7449
rect 6736 7404 6788 7410
rect 6656 7364 6736 7392
rect 7012 7414 7064 7420
rect 7300 7410 7328 7482
rect 6826 7375 6882 7384
rect 7288 7404 7340 7410
rect 6736 7346 6788 7352
rect 7288 7346 7340 7352
rect 6512 7296 6684 7324
rect 6460 7278 6512 7284
rect 6366 7168 6422 7177
rect 6366 7103 6422 7112
rect 6380 7002 6408 7103
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6366 6896 6422 6905
rect 6196 6820 6316 6848
rect 6366 6831 6422 6840
rect 6288 6662 6316 6820
rect 6000 6656 6052 6662
rect 6276 6656 6328 6662
rect 6000 6598 6052 6604
rect 6090 6624 6146 6633
rect 6012 6186 6040 6598
rect 6276 6598 6328 6604
rect 6090 6559 6146 6568
rect 6104 6390 6132 6559
rect 6182 6488 6238 6497
rect 6380 6458 6408 6831
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6182 6423 6238 6432
rect 6368 6452 6420 6458
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 6104 5642 6132 6190
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6104 5302 6132 5578
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 6012 4622 6040 5102
rect 6196 5030 6224 6423
rect 6368 6394 6420 6400
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6288 5574 6316 6326
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 5370 6316 5510
rect 6472 5370 6500 6598
rect 6564 6497 6592 6734
rect 6550 6488 6606 6497
rect 6550 6423 6606 6432
rect 6550 6080 6606 6089
rect 6550 6015 6606 6024
rect 6564 5914 6592 6015
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6380 5030 6408 5170
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6182 4856 6238 4865
rect 6182 4791 6184 4800
rect 6236 4791 6238 4800
rect 6184 4762 6236 4768
rect 6552 4752 6604 4758
rect 6656 4740 6684 7296
rect 6872 7100 7180 7109
rect 6872 7098 6878 7100
rect 6934 7098 6958 7100
rect 7014 7098 7038 7100
rect 7094 7098 7118 7100
rect 7174 7098 7180 7100
rect 6934 7046 6936 7098
rect 7116 7046 7118 7098
rect 6872 7044 6878 7046
rect 6934 7044 6958 7046
rect 7014 7044 7038 7046
rect 7094 7044 7118 7046
rect 7174 7044 7180 7046
rect 6872 7035 7180 7044
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 7012 6996 7064 7002
rect 7300 6984 7328 7346
rect 7012 6938 7064 6944
rect 7208 6956 7328 6984
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6748 6730 6776 6870
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6840 6458 6868 6938
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6932 6497 6960 6734
rect 7024 6730 7052 6938
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6918 6488 6974 6497
rect 6828 6452 6880 6458
rect 6918 6423 6974 6432
rect 6828 6394 6880 6400
rect 6932 6100 6960 6423
rect 7208 6322 7236 6956
rect 7286 6896 7342 6905
rect 7286 6831 7342 6840
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 6118 7236 6258
rect 6748 6072 6960 6100
rect 7196 6112 7248 6118
rect 6748 5710 6776 6072
rect 7196 6054 7248 6060
rect 6872 6012 7180 6021
rect 6872 6010 6878 6012
rect 6934 6010 6958 6012
rect 7014 6010 7038 6012
rect 7094 6010 7118 6012
rect 7174 6010 7180 6012
rect 6934 5958 6936 6010
rect 7116 5958 7118 6010
rect 6872 5956 6878 5958
rect 6934 5956 6958 5958
rect 7014 5956 7038 5958
rect 7094 5956 7118 5958
rect 7174 5956 7180 5958
rect 6872 5947 7180 5956
rect 7300 5778 7328 6831
rect 7392 6100 7420 9590
rect 7484 8974 7512 10474
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 7857 7512 8774
rect 7576 8634 7604 13110
rect 7668 12850 7696 14991
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7760 13814 7788 13874
rect 7760 13786 7880 13814
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7760 12730 7788 13398
rect 7668 12702 7788 12730
rect 7668 12442 7696 12702
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7668 12170 7696 12378
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7668 11082 7696 12106
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7654 10296 7710 10305
rect 7654 10231 7710 10240
rect 7668 10062 7696 10231
rect 7760 10062 7788 12582
rect 7852 12322 7880 13786
rect 7944 12442 7972 15914
rect 8846 15260 9154 15269
rect 8846 15258 8852 15260
rect 8908 15258 8932 15260
rect 8988 15258 9012 15260
rect 9068 15258 9092 15260
rect 9148 15258 9154 15260
rect 8908 15206 8910 15258
rect 9090 15206 9092 15258
rect 8846 15204 8852 15206
rect 8908 15204 8932 15206
rect 8988 15204 9012 15206
rect 9068 15204 9092 15206
rect 9148 15204 9154 15206
rect 8846 15195 9154 15204
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8036 13433 8064 13806
rect 8022 13424 8078 13433
rect 8022 13359 8078 13368
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12918 8064 13126
rect 8024 12912 8076 12918
rect 8024 12854 8076 12860
rect 8114 12880 8170 12889
rect 8114 12815 8170 12824
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 8036 12617 8064 12718
rect 8022 12608 8078 12617
rect 8022 12543 8078 12552
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7852 12294 7972 12322
rect 7944 11801 7972 12294
rect 7930 11792 7986 11801
rect 8036 11762 8064 12543
rect 8128 12238 8156 12815
rect 8220 12374 8248 13874
rect 8312 12986 8340 14758
rect 8404 13326 8432 14826
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8312 12442 8340 12922
rect 8496 12730 8524 15098
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8588 12968 8616 15030
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8680 13297 8708 13874
rect 8772 13394 8800 14894
rect 8846 14172 9154 14181
rect 8846 14170 8852 14172
rect 8908 14170 8932 14172
rect 8988 14170 9012 14172
rect 9068 14170 9092 14172
rect 9148 14170 9154 14172
rect 8908 14118 8910 14170
rect 9090 14118 9092 14170
rect 8846 14116 8852 14118
rect 8908 14116 8932 14118
rect 8988 14116 9012 14118
rect 9068 14116 9092 14118
rect 9148 14116 9154 14118
rect 8846 14107 9154 14116
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8666 13288 8722 13297
rect 8666 13223 8722 13232
rect 8846 13084 9154 13093
rect 8846 13082 8852 13084
rect 8908 13082 8932 13084
rect 8988 13082 9012 13084
rect 9068 13082 9092 13084
rect 9148 13082 9154 13084
rect 8908 13030 8910 13082
rect 9090 13030 9092 13082
rect 8846 13028 8852 13030
rect 8908 13028 8932 13030
rect 8988 13028 9012 13030
rect 9068 13028 9092 13030
rect 9148 13028 9154 13030
rect 8846 13019 9154 13028
rect 8588 12940 8984 12968
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8496 12702 8800 12730
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8116 12096 8168 12102
rect 8220 12084 8248 12310
rect 8220 12056 8340 12084
rect 8116 12038 8168 12044
rect 7930 11727 7986 11736
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7838 11656 7894 11665
rect 7838 11591 7894 11600
rect 7852 11257 7880 11591
rect 7838 11248 7894 11257
rect 7838 11183 7894 11192
rect 8024 11212 8076 11218
rect 7852 11150 7880 11183
rect 8024 11154 8076 11160
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7668 9353 7696 9998
rect 7654 9344 7710 9353
rect 7654 9279 7710 9288
rect 7654 9208 7710 9217
rect 7654 9143 7710 9152
rect 7668 9110 7696 9143
rect 7656 9104 7708 9110
rect 7852 9092 7880 10066
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7944 9178 7972 9386
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7656 9046 7708 9052
rect 7760 9064 7880 9092
rect 8036 9081 8064 11154
rect 8128 10810 8156 12038
rect 8312 11830 8340 12056
rect 8300 11824 8352 11830
rect 8206 11792 8262 11801
rect 8300 11766 8352 11772
rect 8206 11727 8262 11736
rect 8220 11694 8248 11727
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8404 11082 8432 12582
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8300 10668 8352 10674
rect 8404 10656 8432 11018
rect 8352 10628 8432 10656
rect 8300 10610 8352 10616
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8022 9072 8078 9081
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7562 8392 7618 8401
rect 7562 8327 7564 8336
rect 7616 8327 7618 8336
rect 7564 8298 7616 8304
rect 7668 8090 7696 9046
rect 7760 8922 7788 9064
rect 8022 9007 8078 9016
rect 7760 8894 7880 8922
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7656 8084 7708 8090
rect 7576 8044 7656 8072
rect 7470 7848 7526 7857
rect 7470 7783 7526 7792
rect 7484 7342 7512 7783
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7576 6984 7604 8044
rect 7656 8026 7708 8032
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7484 6956 7604 6984
rect 7484 6866 7512 6956
rect 7562 6896 7618 6905
rect 7472 6860 7524 6866
rect 7562 6831 7564 6840
rect 7472 6802 7524 6808
rect 7616 6831 7618 6840
rect 7564 6802 7616 6808
rect 7481 6112 7533 6118
rect 7392 6072 7481 6100
rect 7481 6054 7533 6060
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7380 5704 7432 5710
rect 7576 5681 7604 5782
rect 7380 5646 7432 5652
rect 7562 5672 7618 5681
rect 6932 5370 6960 5646
rect 7392 5574 7420 5646
rect 7562 5607 7618 5616
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7116 5234 7144 5510
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 6748 5098 6776 5170
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6748 4826 6776 5034
rect 6872 4924 7180 4933
rect 6872 4922 6878 4924
rect 6934 4922 6958 4924
rect 7014 4922 7038 4924
rect 7094 4922 7118 4924
rect 7174 4922 7180 4924
rect 6934 4870 6936 4922
rect 7116 4870 7118 4922
rect 6872 4868 6878 4870
rect 6934 4868 6958 4870
rect 7014 4868 7038 4870
rect 7094 4868 7118 4870
rect 7174 4868 7180 4870
rect 6872 4859 7180 4868
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6604 4712 6684 4740
rect 6552 4694 6604 4700
rect 7208 4690 7236 5306
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6184 4616 6236 4622
rect 6644 4616 6696 4622
rect 6184 4558 6236 4564
rect 6642 4584 6644 4593
rect 6696 4584 6698 4593
rect 6012 4214 6040 4558
rect 6000 4208 6052 4214
rect 5722 4176 5778 4185
rect 6000 4150 6052 4156
rect 6196 4146 6224 4558
rect 6642 4519 6698 4528
rect 7300 4185 7328 5034
rect 7286 4176 7342 4185
rect 5722 4111 5778 4120
rect 6184 4140 6236 4146
rect 5630 3904 5686 3913
rect 5630 3839 5686 3848
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4898 3292 5206 3301
rect 4898 3290 4904 3292
rect 4960 3290 4984 3292
rect 5040 3290 5064 3292
rect 5120 3290 5144 3292
rect 5200 3290 5206 3292
rect 4960 3238 4962 3290
rect 5142 3238 5144 3290
rect 4898 3236 4904 3238
rect 4960 3236 4984 3238
rect 5040 3236 5064 3238
rect 5120 3236 5144 3238
rect 5200 3236 5206 3238
rect 4898 3227 5206 3236
rect 5736 2446 5764 4111
rect 7286 4111 7342 4120
rect 6184 4082 6236 4088
rect 7392 3942 7420 5510
rect 7668 5409 7696 7346
rect 7760 6798 7788 8774
rect 7852 8090 7880 8894
rect 8024 8832 8076 8838
rect 7944 8792 8024 8820
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7852 7732 7880 7890
rect 7944 7886 7972 8792
rect 8024 8774 8076 8780
rect 8024 8492 8076 8498
rect 8128 8480 8156 9658
rect 8206 9480 8262 9489
rect 8206 9415 8208 9424
rect 8260 9415 8262 9424
rect 8208 9386 8260 9392
rect 8206 9344 8262 9353
rect 8206 9279 8262 9288
rect 8220 8974 8248 9279
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8220 8809 8248 8910
rect 8206 8800 8262 8809
rect 8206 8735 8262 8744
rect 8076 8452 8248 8480
rect 8024 8434 8076 8440
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7852 7704 7972 7732
rect 7838 7576 7894 7585
rect 7838 7511 7894 7520
rect 7852 7177 7880 7511
rect 7838 7168 7894 7177
rect 7838 7103 7894 7112
rect 7944 6882 7972 7704
rect 7852 6854 7972 6882
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7760 5710 7788 6326
rect 7852 6186 7880 6854
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7748 5704 7800 5710
rect 7840 5704 7892 5710
rect 7748 5646 7800 5652
rect 7838 5672 7840 5681
rect 7892 5672 7894 5681
rect 7654 5400 7710 5409
rect 7654 5335 7710 5344
rect 7760 4282 7788 5646
rect 7838 5607 7894 5616
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 6872 3836 7180 3845
rect 6872 3834 6878 3836
rect 6934 3834 6958 3836
rect 7014 3834 7038 3836
rect 7094 3834 7118 3836
rect 7174 3834 7180 3836
rect 6934 3782 6936 3834
rect 7116 3782 7118 3834
rect 6872 3780 6878 3782
rect 6934 3780 6958 3782
rect 7014 3780 7038 3782
rect 7094 3780 7118 3782
rect 7174 3780 7180 3782
rect 6872 3771 7180 3780
rect 7944 3058 7972 6734
rect 8036 5574 8064 8298
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8128 6730 8156 7958
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8128 6322 8156 6666
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8128 5166 8156 6054
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8220 5030 8248 8452
rect 8312 8090 8340 9998
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8404 7886 8432 9862
rect 8496 9042 8524 12582
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8588 12073 8616 12106
rect 8574 12064 8630 12073
rect 8574 11999 8630 12008
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8588 9518 8616 11834
rect 8680 10198 8708 12106
rect 8772 11642 8800 12702
rect 8864 12481 8892 12786
rect 8956 12714 8984 12940
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 9048 12753 9076 12854
rect 9034 12744 9090 12753
rect 8944 12708 8996 12714
rect 9034 12679 9090 12688
rect 8944 12650 8996 12656
rect 8850 12472 8906 12481
rect 8850 12407 8906 12416
rect 8956 12238 8984 12650
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9048 12170 9076 12679
rect 9232 12646 9260 16594
rect 10820 15804 11128 15813
rect 10820 15802 10826 15804
rect 10882 15802 10906 15804
rect 10962 15802 10986 15804
rect 11042 15802 11066 15804
rect 11122 15802 11128 15804
rect 10882 15750 10884 15802
rect 11064 15750 11066 15802
rect 10820 15748 10826 15750
rect 10882 15748 10906 15750
rect 10962 15748 10986 15750
rect 11042 15748 11066 15750
rect 11122 15748 11128 15750
rect 10820 15739 11128 15748
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9126 12336 9182 12345
rect 9324 12322 9352 14418
rect 9600 13530 9628 15642
rect 10820 14716 11128 14725
rect 10820 14714 10826 14716
rect 10882 14714 10906 14716
rect 10962 14714 10986 14716
rect 11042 14714 11066 14716
rect 11122 14714 11128 14716
rect 10882 14662 10884 14714
rect 11064 14662 11066 14714
rect 10820 14660 10826 14662
rect 10882 14660 10906 14662
rect 10962 14660 10986 14662
rect 11042 14660 11066 14662
rect 11122 14660 11128 14662
rect 10820 14651 11128 14660
rect 10598 14376 10654 14385
rect 10598 14311 10654 14320
rect 10322 13968 10378 13977
rect 10322 13903 10378 13912
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9508 12481 9536 12582
rect 9494 12472 9550 12481
rect 9494 12407 9550 12416
rect 9692 12345 9720 12718
rect 9678 12336 9734 12345
rect 9324 12294 9536 12322
rect 9126 12271 9182 12280
rect 9140 12238 9168 12271
rect 9128 12232 9180 12238
rect 9404 12232 9456 12238
rect 9180 12192 9352 12220
rect 9128 12174 9180 12180
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 8846 11996 9154 12005
rect 8846 11994 8852 11996
rect 8908 11994 8932 11996
rect 8988 11994 9012 11996
rect 9068 11994 9092 11996
rect 9148 11994 9154 11996
rect 8908 11942 8910 11994
rect 9090 11942 9092 11994
rect 8846 11940 8852 11942
rect 8908 11940 8932 11942
rect 8988 11940 9012 11942
rect 9068 11940 9092 11942
rect 9148 11940 9154 11942
rect 8846 11931 9154 11940
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 8944 11688 8996 11694
rect 8772 11614 8892 11642
rect 8944 11630 8996 11636
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8772 10713 8800 11494
rect 8864 11257 8892 11614
rect 8956 11558 8984 11630
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8850 11248 8906 11257
rect 8850 11183 8906 11192
rect 9048 11121 9076 11698
rect 9324 11642 9352 12192
rect 9404 12174 9456 12180
rect 9508 12186 9536 12294
rect 9678 12271 9734 12280
rect 9416 11880 9444 12174
rect 9508 12158 9720 12186
rect 9692 12102 9720 12158
rect 9680 12096 9732 12102
rect 9586 12064 9642 12073
rect 9680 12038 9732 12044
rect 9586 11999 9642 12008
rect 9416 11852 9536 11880
rect 9402 11792 9458 11801
rect 9402 11727 9404 11736
rect 9456 11727 9458 11736
rect 9404 11698 9456 11704
rect 9232 11614 9352 11642
rect 9126 11520 9182 11529
rect 9126 11455 9182 11464
rect 9140 11218 9168 11455
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9232 11121 9260 11614
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9034 11112 9090 11121
rect 9034 11047 9090 11056
rect 9218 11112 9274 11121
rect 9218 11047 9274 11056
rect 8846 10908 9154 10917
rect 8846 10906 8852 10908
rect 8908 10906 8932 10908
rect 8988 10906 9012 10908
rect 9068 10906 9092 10908
rect 9148 10906 9154 10908
rect 8908 10854 8910 10906
rect 9090 10854 9092 10906
rect 8846 10852 8852 10854
rect 8908 10852 8932 10854
rect 8988 10852 9012 10854
rect 9068 10852 9092 10854
rect 9148 10852 9154 10854
rect 8846 10843 9154 10852
rect 8758 10704 8814 10713
rect 8758 10639 8814 10648
rect 8942 10704 8998 10713
rect 8942 10639 8998 10648
rect 8956 10305 8984 10639
rect 8942 10296 8998 10305
rect 8942 10231 8998 10240
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8680 9586 8708 10134
rect 9232 9874 9260 11047
rect 9324 10742 9352 11494
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9508 10282 9536 11852
rect 9600 11150 9628 11999
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9678 11520 9734 11529
rect 9678 11455 9734 11464
rect 9692 11218 9720 11455
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9416 10254 9536 10282
rect 9416 10198 9444 10254
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9232 9846 9352 9874
rect 8846 9820 9154 9829
rect 8846 9818 8852 9820
rect 8908 9818 8932 9820
rect 8988 9818 9012 9820
rect 9068 9818 9092 9820
rect 9148 9818 9154 9820
rect 8908 9766 8910 9818
rect 9090 9766 9092 9818
rect 8846 9764 8852 9766
rect 8908 9764 8932 9766
rect 8988 9764 9012 9766
rect 9068 9764 9092 9766
rect 9148 9764 9154 9766
rect 8846 9755 9154 9764
rect 9324 9602 9352 9846
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 9048 9574 9352 9602
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8574 9344 8630 9353
rect 8574 9279 8630 9288
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8588 8974 8616 9279
rect 8666 9072 8722 9081
rect 8666 9007 8722 9016
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8496 8566 8524 8774
rect 8574 8664 8630 8673
rect 8574 8599 8630 8608
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8390 7712 8446 7721
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8312 3534 8340 7686
rect 8390 7647 8446 7656
rect 8404 7478 8432 7647
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8404 6202 8432 6734
rect 8496 6361 8524 7958
rect 8482 6352 8538 6361
rect 8588 6322 8616 8599
rect 8680 8498 8708 9007
rect 9048 8906 9076 9574
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9220 9512 9272 9518
rect 9416 9500 9444 10134
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9272 9472 9444 9500
rect 9220 9454 9272 9460
rect 9140 9058 9168 9454
rect 9404 9376 9456 9382
rect 9402 9344 9404 9353
rect 9456 9344 9458 9353
rect 9402 9279 9458 9288
rect 9140 9030 9444 9058
rect 9128 8968 9180 8974
rect 9180 8916 9352 8922
rect 9128 8910 9352 8916
rect 9036 8900 9088 8906
rect 9140 8894 9352 8910
rect 9036 8842 9088 8848
rect 9324 8838 9352 8894
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 8846 8732 9154 8741
rect 8846 8730 8852 8732
rect 8908 8730 8932 8732
rect 8988 8730 9012 8732
rect 9068 8730 9092 8732
rect 9148 8730 9154 8732
rect 8908 8678 8910 8730
rect 9090 8678 9092 8730
rect 8846 8676 8852 8678
rect 8908 8676 8932 8678
rect 8988 8676 9012 8678
rect 9068 8676 9092 8678
rect 9148 8676 9154 8678
rect 8846 8667 9154 8676
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8680 6866 8708 8298
rect 8772 7546 8800 8298
rect 8956 8129 8984 8434
rect 9048 8401 9076 8502
rect 9034 8392 9090 8401
rect 9034 8327 9090 8336
rect 8942 8120 8998 8129
rect 8942 8055 8998 8064
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 8846 7644 9154 7653
rect 8846 7642 8852 7644
rect 8908 7642 8932 7644
rect 8988 7642 9012 7644
rect 9068 7642 9092 7644
rect 9148 7642 9154 7644
rect 8908 7590 8910 7642
rect 9090 7590 9092 7642
rect 8846 7588 8852 7590
rect 8908 7588 8932 7590
rect 8988 7588 9012 7590
rect 9068 7588 9092 7590
rect 9148 7588 9154 7590
rect 8846 7579 9154 7588
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 9034 7440 9090 7449
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8772 7002 8800 7346
rect 8956 7342 8984 7414
rect 9034 7375 9090 7384
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 9048 7002 9076 7375
rect 9128 7268 9180 7274
rect 9232 7256 9260 7958
rect 9180 7228 9260 7256
rect 9128 7210 9180 7216
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8482 6287 8538 6296
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8680 6254 8708 6802
rect 8772 6361 8800 6938
rect 9324 6934 9352 8774
rect 9416 8090 9444 9030
rect 9508 8974 9536 10066
rect 9600 10010 9628 11086
rect 9678 10840 9734 10849
rect 9784 10810 9812 11630
rect 9876 11354 9904 13262
rect 9968 11354 9996 13806
rect 10138 12880 10194 12889
rect 10048 12844 10100 12850
rect 10138 12815 10194 12824
rect 10048 12786 10100 12792
rect 10060 12238 10088 12786
rect 10152 12646 10180 12815
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 10060 11286 10088 12174
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10152 11898 10180 12038
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10152 11665 10180 11698
rect 10244 11694 10272 12582
rect 10232 11688 10284 11694
rect 10138 11656 10194 11665
rect 10232 11630 10284 11636
rect 10138 11591 10194 11600
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10138 11248 10194 11257
rect 10244 11234 10272 11630
rect 10336 11354 10364 13903
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10244 11206 10364 11234
rect 10138 11183 10194 11192
rect 10152 11132 10180 11183
rect 10232 11144 10284 11150
rect 10152 11104 10232 11132
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9678 10775 9680 10784
rect 9732 10775 9734 10784
rect 9772 10804 9824 10810
rect 9680 10746 9732 10752
rect 9772 10746 9824 10752
rect 9876 10441 9904 10950
rect 10048 10464 10100 10470
rect 9862 10432 9918 10441
rect 10048 10406 10100 10412
rect 9862 10367 9918 10376
rect 9864 10056 9916 10062
rect 9600 9982 9812 10010
rect 9864 9998 9916 10004
rect 9680 9920 9732 9926
rect 9586 9888 9642 9897
rect 9680 9862 9732 9868
rect 9586 9823 9642 9832
rect 9600 9722 9628 9823
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9692 9217 9720 9862
rect 9678 9208 9734 9217
rect 9784 9178 9812 9982
rect 9876 9654 9904 9998
rect 10060 9761 10088 10406
rect 10046 9752 10102 9761
rect 9956 9716 10008 9722
rect 10046 9687 10102 9696
rect 9956 9658 10008 9664
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9678 9143 9734 9152
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9508 8634 9536 8910
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9600 8514 9628 9046
rect 9784 8634 9812 9114
rect 9876 9081 9904 9590
rect 9968 9489 9996 9658
rect 9954 9480 10010 9489
rect 9954 9415 10010 9424
rect 10152 9353 10180 11104
rect 10232 11086 10284 11092
rect 10336 10674 10364 11206
rect 10324 10668 10376 10674
rect 10428 10658 10456 12378
rect 10520 12170 10548 13194
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10506 11520 10562 11529
rect 10506 11455 10562 11464
rect 10520 11286 10548 11455
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10612 11150 10640 14311
rect 10820 13628 11128 13637
rect 10820 13626 10826 13628
rect 10882 13626 10906 13628
rect 10962 13626 10986 13628
rect 11042 13626 11066 13628
rect 11122 13626 11128 13628
rect 10882 13574 10884 13626
rect 11064 13574 11066 13626
rect 10820 13572 10826 13574
rect 10882 13572 10906 13574
rect 10962 13572 10986 13574
rect 11042 13572 11066 13574
rect 11122 13572 11128 13574
rect 10820 13563 11128 13572
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10704 12306 10732 13330
rect 11072 12850 11100 13466
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11256 12646 11284 13126
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 10820 12540 11128 12549
rect 10820 12538 10826 12540
rect 10882 12538 10906 12540
rect 10962 12538 10986 12540
rect 11042 12538 11066 12540
rect 11122 12538 11128 12540
rect 10882 12486 10884 12538
rect 11064 12486 11066 12538
rect 10820 12484 10826 12486
rect 10882 12484 10906 12486
rect 10962 12484 10986 12486
rect 11042 12484 11066 12486
rect 11122 12484 11128 12486
rect 10820 12475 11128 12484
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10796 12345 10824 12378
rect 10782 12336 10838 12345
rect 10692 12300 10744 12306
rect 10782 12271 10838 12280
rect 10692 12242 10744 12248
rect 10704 11801 10732 12242
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10690 11792 10746 11801
rect 10690 11727 10746 11736
rect 10796 11676 10824 12106
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10704 11648 10824 11676
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10704 10996 10732 11648
rect 10820 11452 11128 11461
rect 10820 11450 10826 11452
rect 10882 11450 10906 11452
rect 10962 11450 10986 11452
rect 11042 11450 11066 11452
rect 11122 11450 11128 11452
rect 10882 11398 10884 11450
rect 11064 11398 11066 11450
rect 10820 11396 10826 11398
rect 10882 11396 10906 11398
rect 10962 11396 10986 11398
rect 11042 11396 11066 11398
rect 11122 11396 11128 11398
rect 10820 11387 11128 11396
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10796 11121 10824 11290
rect 11164 11257 11192 12038
rect 11150 11248 11206 11257
rect 11150 11183 11206 11192
rect 11164 11150 11192 11183
rect 11152 11144 11204 11150
rect 10782 11112 10838 11121
rect 11152 11086 11204 11092
rect 10782 11047 10784 11056
rect 10836 11047 10838 11056
rect 10784 11018 10836 11024
rect 10520 10968 10732 10996
rect 10796 10987 10824 11018
rect 11256 11014 11284 12582
rect 11348 12442 11376 17206
rect 14768 16892 15076 16901
rect 14768 16890 14774 16892
rect 14830 16890 14854 16892
rect 14910 16890 14934 16892
rect 14990 16890 15014 16892
rect 15070 16890 15076 16892
rect 14830 16838 14832 16890
rect 15012 16838 15014 16890
rect 14768 16836 14774 16838
rect 14830 16836 14854 16838
rect 14910 16836 14934 16838
rect 14990 16836 15014 16838
rect 15070 16836 15076 16838
rect 14768 16827 15076 16836
rect 12794 16348 13102 16357
rect 12794 16346 12800 16348
rect 12856 16346 12880 16348
rect 12936 16346 12960 16348
rect 13016 16346 13040 16348
rect 13096 16346 13102 16348
rect 12856 16294 12858 16346
rect 13038 16294 13040 16346
rect 12794 16292 12800 16294
rect 12856 16292 12880 16294
rect 12936 16292 12960 16294
rect 13016 16292 13040 16294
rect 13096 16292 13102 16294
rect 12794 16283 13102 16292
rect 14768 15804 15076 15813
rect 14768 15802 14774 15804
rect 14830 15802 14854 15804
rect 14910 15802 14934 15804
rect 14990 15802 15014 15804
rect 15070 15802 15076 15804
rect 14830 15750 14832 15802
rect 15012 15750 15014 15802
rect 14768 15748 14774 15750
rect 14830 15748 14854 15750
rect 14910 15748 14934 15750
rect 14990 15748 15014 15750
rect 15070 15748 15076 15750
rect 14768 15739 15076 15748
rect 12794 15260 13102 15269
rect 12794 15258 12800 15260
rect 12856 15258 12880 15260
rect 12936 15258 12960 15260
rect 13016 15258 13040 15260
rect 13096 15258 13102 15260
rect 12856 15206 12858 15258
rect 13038 15206 13040 15258
rect 12794 15204 12800 15206
rect 12856 15204 12880 15206
rect 12936 15204 12960 15206
rect 13016 15204 13040 15206
rect 13096 15204 13102 15206
rect 12794 15195 13102 15204
rect 14768 14716 15076 14725
rect 14768 14714 14774 14716
rect 14830 14714 14854 14716
rect 14910 14714 14934 14716
rect 14990 14714 15014 14716
rect 15070 14714 15076 14716
rect 14830 14662 14832 14714
rect 15012 14662 15014 14714
rect 14768 14660 14774 14662
rect 14830 14660 14854 14662
rect 14910 14660 14934 14662
rect 14990 14660 15014 14662
rect 15070 14660 15076 14662
rect 14768 14651 15076 14660
rect 12794 14172 13102 14181
rect 12794 14170 12800 14172
rect 12856 14170 12880 14172
rect 12936 14170 12960 14172
rect 13016 14170 13040 14172
rect 13096 14170 13102 14172
rect 12856 14118 12858 14170
rect 13038 14118 13040 14170
rect 12794 14116 12800 14118
rect 12856 14116 12880 14118
rect 12936 14116 12960 14118
rect 13016 14116 13040 14118
rect 13096 14116 13102 14118
rect 12794 14107 13102 14116
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 10876 11008 10928 11014
rect 10324 10610 10376 10616
rect 10416 10652 10468 10658
rect 10232 10600 10284 10606
rect 10416 10594 10468 10600
rect 10232 10542 10284 10548
rect 10244 9722 10272 10542
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10520 10010 10548 10968
rect 10876 10950 10928 10956
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 10888 10849 10916 10950
rect 10874 10840 10930 10849
rect 10874 10775 10930 10784
rect 11256 10742 11284 10950
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 10796 10452 10824 10678
rect 11150 10568 11206 10577
rect 11150 10503 11206 10512
rect 10612 10424 10824 10452
rect 10612 10266 10640 10424
rect 10820 10364 11128 10373
rect 10820 10362 10826 10364
rect 10882 10362 10906 10364
rect 10962 10362 10986 10364
rect 11042 10362 11066 10364
rect 11122 10362 11128 10364
rect 10882 10310 10884 10362
rect 11064 10310 11066 10362
rect 10820 10308 10826 10310
rect 10882 10308 10906 10310
rect 10962 10308 10986 10310
rect 11042 10308 11066 10310
rect 11122 10308 11128 10310
rect 10690 10296 10746 10305
rect 10820 10299 11128 10308
rect 10600 10260 10652 10266
rect 10690 10231 10746 10240
rect 10600 10202 10652 10208
rect 10704 10146 10732 10231
rect 10704 10118 10824 10146
rect 10796 10062 10824 10118
rect 10784 10056 10836 10062
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10138 9344 10194 9353
rect 9968 9302 10138 9330
rect 9862 9072 9918 9081
rect 9862 9007 9918 9016
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9496 8492 9548 8498
rect 9600 8486 9720 8514
rect 9496 8434 9548 8440
rect 9508 8294 9536 8434
rect 9692 8344 9720 8486
rect 9772 8492 9824 8498
rect 9968 8480 9996 9302
rect 10138 9279 10194 9288
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9824 8452 9996 8480
rect 9772 8434 9824 8440
rect 9600 8316 9720 8344
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9416 7313 9444 7754
rect 9402 7304 9458 7313
rect 9402 7239 9458 7248
rect 9404 7200 9456 7206
rect 9402 7168 9404 7177
rect 9456 7168 9458 7177
rect 9402 7103 9458 7112
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 8846 6556 9154 6565
rect 8846 6554 8852 6556
rect 8908 6554 8932 6556
rect 8988 6554 9012 6556
rect 9068 6554 9092 6556
rect 9148 6554 9154 6556
rect 8908 6502 8910 6554
rect 9090 6502 9092 6554
rect 8846 6500 8852 6502
rect 8908 6500 8932 6502
rect 8988 6500 9012 6502
rect 9068 6500 9092 6502
rect 9148 6500 9154 6502
rect 8846 6491 9154 6500
rect 9232 6390 9260 6734
rect 9220 6384 9272 6390
rect 8758 6352 8814 6361
rect 9220 6326 9272 6332
rect 8758 6287 8814 6296
rect 8668 6248 8720 6254
rect 8404 6174 8524 6202
rect 8668 6190 8720 6196
rect 8758 6216 8814 6225
rect 8496 5778 8524 6174
rect 8758 6151 8760 6160
rect 8812 6151 8814 6160
rect 8760 6122 8812 6128
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8496 5574 8524 5714
rect 8484 5568 8536 5574
rect 8404 5528 8484 5556
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8404 2990 8432 5528
rect 8484 5510 8536 5516
rect 8846 5468 9154 5477
rect 8846 5466 8852 5468
rect 8908 5466 8932 5468
rect 8988 5466 9012 5468
rect 9068 5466 9092 5468
rect 9148 5466 9154 5468
rect 8908 5414 8910 5466
rect 9090 5414 9092 5466
rect 8846 5412 8852 5414
rect 8908 5412 8932 5414
rect 8988 5412 9012 5414
rect 9068 5412 9092 5414
rect 9148 5412 9154 5414
rect 8482 5400 8538 5409
rect 8846 5403 9154 5412
rect 8482 5335 8538 5344
rect 8496 5302 8524 5335
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 9508 4758 9536 8230
rect 9600 7002 9628 8316
rect 9876 7886 9904 8452
rect 10060 8401 10088 8774
rect 10046 8392 10102 8401
rect 10046 8327 10102 8336
rect 9864 7880 9916 7886
rect 9916 7840 9996 7868
rect 9864 7822 9916 7828
rect 9864 7744 9916 7750
rect 9678 7712 9734 7721
rect 9864 7686 9916 7692
rect 9678 7647 9734 7656
rect 9692 7478 9720 7647
rect 9876 7585 9904 7686
rect 9862 7576 9918 7585
rect 9862 7511 9918 7520
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9784 6882 9812 7346
rect 9692 6854 9812 6882
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9600 6254 9628 6734
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9692 5778 9720 6854
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 8846 4380 9154 4389
rect 8846 4378 8852 4380
rect 8908 4378 8932 4380
rect 8988 4378 9012 4380
rect 9068 4378 9092 4380
rect 9148 4378 9154 4380
rect 8908 4326 8910 4378
rect 9090 4326 9092 4378
rect 8846 4324 8852 4326
rect 8908 4324 8932 4326
rect 8988 4324 9012 4326
rect 9068 4324 9092 4326
rect 9148 4324 9154 4326
rect 8846 4315 9154 4324
rect 8846 3292 9154 3301
rect 8846 3290 8852 3292
rect 8908 3290 8932 3292
rect 8988 3290 9012 3292
rect 9068 3290 9092 3292
rect 9148 3290 9154 3292
rect 8908 3238 8910 3290
rect 9090 3238 9092 3290
rect 8846 3236 8852 3238
rect 8908 3236 8932 3238
rect 8988 3236 9012 3238
rect 9068 3236 9092 3238
rect 9148 3236 9154 3238
rect 8846 3227 9154 3236
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 9784 2854 9812 6734
rect 9876 4486 9904 7511
rect 9968 6662 9996 7840
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 10060 6390 10088 7346
rect 10152 6866 10180 9114
rect 10244 7546 10272 9658
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10336 6905 10364 9998
rect 10428 9674 10456 9998
rect 10520 9982 10732 10010
rect 10784 9998 10836 10004
rect 10428 9646 10640 9674
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 9217 10548 9522
rect 10612 9518 10640 9646
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10506 9208 10562 9217
rect 10506 9143 10508 9152
rect 10560 9143 10562 9152
rect 10508 9114 10560 9120
rect 10520 9083 10548 9114
rect 10612 9110 10640 9454
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10704 9058 10732 9982
rect 10820 9276 11128 9285
rect 10820 9274 10826 9276
rect 10882 9274 10906 9276
rect 10962 9274 10986 9276
rect 11042 9274 11066 9276
rect 11122 9274 11128 9276
rect 10882 9222 10884 9274
rect 11064 9222 11066 9274
rect 10820 9220 10826 9222
rect 10882 9220 10906 9222
rect 10962 9220 10986 9222
rect 11042 9220 11066 9222
rect 11122 9220 11128 9222
rect 10820 9211 11128 9220
rect 11164 9178 11192 10503
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 10704 9030 11008 9058
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10428 8430 10456 8842
rect 10508 8832 10560 8838
rect 10612 8809 10640 8910
rect 10508 8774 10560 8780
rect 10598 8800 10654 8809
rect 10520 8634 10548 8774
rect 10598 8735 10654 8744
rect 10782 8800 10838 8809
rect 10782 8735 10838 8744
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10414 8256 10470 8265
rect 10414 8191 10470 8200
rect 10428 7546 10456 8191
rect 10520 7886 10548 8298
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10612 7410 10640 7822
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10322 6896 10378 6905
rect 10140 6860 10192 6866
rect 10322 6831 10378 6840
rect 10140 6802 10192 6808
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 10520 5710 10548 7346
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10612 5642 10640 7346
rect 10704 6458 10732 8434
rect 10796 8294 10824 8735
rect 10874 8664 10930 8673
rect 10874 8599 10930 8608
rect 10888 8498 10916 8599
rect 10980 8566 11008 9030
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11072 8945 11100 8978
rect 11256 8945 11284 9590
rect 11348 9450 11376 11698
rect 11440 10656 11468 12786
rect 11624 12434 11652 13874
rect 14768 13628 15076 13637
rect 14768 13626 14774 13628
rect 14830 13626 14854 13628
rect 14910 13626 14934 13628
rect 14990 13626 15014 13628
rect 15070 13626 15076 13628
rect 14830 13574 14832 13626
rect 15012 13574 15014 13626
rect 14768 13572 14774 13574
rect 14830 13572 14854 13574
rect 14910 13572 14934 13574
rect 14990 13572 15014 13574
rect 15070 13572 15076 13574
rect 14768 13563 15076 13572
rect 12794 13084 13102 13093
rect 12794 13082 12800 13084
rect 12856 13082 12880 13084
rect 12936 13082 12960 13084
rect 13016 13082 13040 13084
rect 13096 13082 13102 13084
rect 12856 13030 12858 13082
rect 13038 13030 13040 13082
rect 12794 13028 12800 13030
rect 12856 13028 12880 13030
rect 12936 13028 12960 13030
rect 13016 13028 13040 13030
rect 13096 13028 13102 13030
rect 12794 13019 13102 13028
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11624 12406 11928 12434
rect 11520 12232 11572 12238
rect 11518 12200 11520 12209
rect 11572 12200 11574 12209
rect 11518 12135 11574 12144
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11624 11354 11652 11562
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11716 10849 11744 11698
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11702 10840 11758 10849
rect 11702 10775 11758 10784
rect 11440 10628 11560 10656
rect 11532 10554 11560 10628
rect 11428 10532 11480 10538
rect 11532 10526 11652 10554
rect 11428 10474 11480 10480
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11336 8968 11388 8974
rect 11058 8936 11114 8945
rect 11242 8936 11298 8945
rect 11058 8871 11114 8880
rect 11152 8900 11204 8906
rect 11440 8956 11468 10474
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11388 8928 11468 8956
rect 11336 8910 11388 8916
rect 11242 8871 11298 8880
rect 11152 8842 11204 8848
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11072 8294 11100 8774
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10820 8188 11128 8197
rect 10820 8186 10826 8188
rect 10882 8186 10906 8188
rect 10962 8186 10986 8188
rect 11042 8186 11066 8188
rect 11122 8186 11128 8188
rect 10882 8134 10884 8186
rect 11064 8134 11066 8186
rect 10820 8132 10826 8134
rect 10882 8132 10906 8134
rect 10962 8132 10986 8134
rect 11042 8132 11066 8134
rect 11122 8132 11128 8134
rect 10820 8123 11128 8132
rect 11164 7886 11192 8842
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11256 8401 11284 8774
rect 11242 8392 11298 8401
rect 11242 8327 11298 8336
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 10968 7880 11020 7886
rect 11152 7880 11204 7886
rect 11020 7828 11100 7834
rect 10968 7822 11100 7828
rect 11152 7822 11204 7828
rect 10980 7806 11100 7822
rect 11072 7750 11100 7806
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10820 7100 11128 7109
rect 10820 7098 10826 7100
rect 10882 7098 10906 7100
rect 10962 7098 10986 7100
rect 11042 7098 11066 7100
rect 11122 7098 11128 7100
rect 10882 7046 10884 7098
rect 11064 7046 11066 7098
rect 10820 7044 10826 7046
rect 10882 7044 10906 7046
rect 10962 7044 10986 7046
rect 11042 7044 11066 7046
rect 11122 7044 11128 7046
rect 10820 7035 11128 7044
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 11164 6118 11192 7822
rect 11256 7750 11284 8230
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 10820 6012 11128 6021
rect 10820 6010 10826 6012
rect 10882 6010 10906 6012
rect 10962 6010 10986 6012
rect 11042 6010 11066 6012
rect 11122 6010 11128 6012
rect 10882 5958 10884 6010
rect 11064 5958 11066 6010
rect 10820 5956 10826 5958
rect 10882 5956 10906 5958
rect 10962 5956 10986 5958
rect 11042 5956 11066 5958
rect 11122 5956 11128 5958
rect 10820 5947 11128 5956
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10820 4924 11128 4933
rect 10820 4922 10826 4924
rect 10882 4922 10906 4924
rect 10962 4922 10986 4924
rect 11042 4922 11066 4924
rect 11122 4922 11128 4924
rect 10882 4870 10884 4922
rect 11064 4870 11066 4922
rect 10820 4868 10826 4870
rect 10882 4868 10906 4870
rect 10962 4868 10986 4870
rect 11042 4868 11066 4870
rect 11122 4868 11128 4870
rect 10820 4859 11128 4868
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 10820 3836 11128 3845
rect 10820 3834 10826 3836
rect 10882 3834 10906 3836
rect 10962 3834 10986 3836
rect 11042 3834 11066 3836
rect 11122 3834 11128 3836
rect 10882 3782 10884 3834
rect 11064 3782 11066 3834
rect 10820 3780 10826 3782
rect 10882 3780 10906 3782
rect 10962 3780 10986 3782
rect 11042 3780 11066 3782
rect 11122 3780 11128 3782
rect 10820 3771 11128 3780
rect 11256 3738 11284 7686
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11348 3466 11376 8910
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11440 6798 11468 8502
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11532 5234 11560 10202
rect 11624 9518 11652 10526
rect 11808 9897 11836 11494
rect 11900 10266 11928 12406
rect 11992 12238 12020 12922
rect 12254 12744 12310 12753
rect 12164 12708 12216 12714
rect 12254 12679 12310 12688
rect 12164 12650 12216 12656
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12084 12442 12112 12582
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12176 12238 12204 12650
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11886 10024 11942 10033
rect 11886 9959 11942 9968
rect 11794 9888 11850 9897
rect 11794 9823 11850 9832
rect 11612 9512 11664 9518
rect 11664 9460 11744 9466
rect 11612 9454 11744 9460
rect 11624 9438 11744 9454
rect 11716 8838 11744 9438
rect 11794 9072 11850 9081
rect 11794 9007 11850 9016
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11624 7478 11652 8434
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11716 6361 11744 8774
rect 11808 8634 11836 9007
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11900 8090 11928 9959
rect 11992 9081 12020 12174
rect 12072 11008 12124 11014
rect 12070 10976 12072 10985
rect 12124 10976 12126 10985
rect 12070 10911 12126 10920
rect 12176 10810 12204 12174
rect 12268 11150 12296 12679
rect 14768 12540 15076 12549
rect 14768 12538 14774 12540
rect 14830 12538 14854 12540
rect 14910 12538 14934 12540
rect 14990 12538 15014 12540
rect 15070 12538 15076 12540
rect 14830 12486 14832 12538
rect 15012 12486 15014 12538
rect 14768 12484 14774 12486
rect 14830 12484 14854 12486
rect 14910 12484 14934 12486
rect 14990 12484 15014 12486
rect 15070 12484 15076 12486
rect 14768 12475 15076 12484
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12360 11762 12388 12310
rect 12794 11996 13102 12005
rect 12794 11994 12800 11996
rect 12856 11994 12880 11996
rect 12936 11994 12960 11996
rect 13016 11994 13040 11996
rect 13096 11994 13102 11996
rect 12856 11942 12858 11994
rect 13038 11942 13040 11994
rect 12794 11940 12800 11942
rect 12856 11940 12880 11942
rect 12936 11940 12960 11942
rect 13016 11940 13040 11942
rect 13096 11940 13102 11942
rect 12794 11931 13102 11940
rect 13910 11792 13966 11801
rect 12348 11756 12400 11762
rect 13910 11727 13966 11736
rect 12348 11698 12400 11704
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12360 10742 12388 11698
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12438 11248 12494 11257
rect 12438 11183 12494 11192
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12084 10606 12112 10678
rect 12452 10674 12480 11183
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 12268 10470 12296 10610
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12084 9722 12112 9998
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 11978 9072 12034 9081
rect 12084 9042 12112 9386
rect 11978 9007 12034 9016
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11702 6352 11758 6361
rect 11702 6287 11758 6296
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11808 5098 11836 7822
rect 11992 5370 12020 8910
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12176 8537 12204 8570
rect 12162 8528 12218 8537
rect 12162 8463 12218 8472
rect 12268 7274 12296 10134
rect 12452 9722 12480 10610
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12346 9616 12402 9625
rect 12346 9551 12348 9560
rect 12400 9551 12402 9560
rect 12440 9580 12492 9586
rect 12348 9522 12400 9528
rect 12440 9522 12492 9528
rect 12360 8616 12388 9522
rect 12452 9489 12480 9522
rect 12438 9480 12494 9489
rect 12438 9415 12494 9424
rect 12360 8588 12480 8616
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12360 7342 12388 8434
rect 12452 8362 12480 8588
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11796 5092 11848 5098
rect 11796 5034 11848 5040
rect 12452 4554 12480 7890
rect 12544 7313 12572 11018
rect 12636 10062 12664 11290
rect 12716 11144 12768 11150
rect 13544 11144 13596 11150
rect 12716 11086 12768 11092
rect 13450 11112 13506 11121
rect 12728 10674 12756 11086
rect 13360 11076 13412 11082
rect 13544 11086 13596 11092
rect 13450 11047 13506 11056
rect 13360 11018 13412 11024
rect 12794 10908 13102 10917
rect 12794 10906 12800 10908
rect 12856 10906 12880 10908
rect 12936 10906 12960 10908
rect 13016 10906 13040 10908
rect 13096 10906 13102 10908
rect 12856 10854 12858 10906
rect 13038 10854 13040 10906
rect 12794 10852 12800 10854
rect 12856 10852 12880 10854
rect 12936 10852 12960 10854
rect 13016 10852 13040 10854
rect 13096 10852 13102 10854
rect 12794 10843 13102 10852
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10062 12756 10406
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12636 9110 12664 9522
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12636 7954 12664 8910
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12530 7304 12586 7313
rect 12530 7239 12586 7248
rect 12728 6769 12756 9862
rect 12794 9820 13102 9829
rect 12794 9818 12800 9820
rect 12856 9818 12880 9820
rect 12936 9818 12960 9820
rect 13016 9818 13040 9820
rect 13096 9818 13102 9820
rect 12856 9766 12858 9818
rect 13038 9766 13040 9818
rect 12794 9764 12800 9766
rect 12856 9764 12880 9766
rect 12936 9764 12960 9766
rect 13016 9764 13040 9766
rect 13096 9764 13102 9766
rect 12794 9755 13102 9764
rect 12794 8732 13102 8741
rect 12794 8730 12800 8732
rect 12856 8730 12880 8732
rect 12936 8730 12960 8732
rect 13016 8730 13040 8732
rect 13096 8730 13102 8732
rect 12856 8678 12858 8730
rect 13038 8678 13040 8730
rect 12794 8676 12800 8678
rect 12856 8676 12880 8678
rect 12936 8676 12960 8678
rect 13016 8676 13040 8678
rect 13096 8676 13102 8678
rect 12794 8667 13102 8676
rect 13188 8022 13216 10610
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13280 10130 13308 10542
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13280 9586 13308 10066
rect 13372 9654 13400 11018
rect 13464 9722 13492 11047
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13176 8016 13228 8022
rect 13556 7993 13584 11086
rect 13924 10742 13952 11727
rect 14768 11452 15076 11461
rect 14768 11450 14774 11452
rect 14830 11450 14854 11452
rect 14910 11450 14934 11452
rect 14990 11450 15014 11452
rect 15070 11450 15076 11452
rect 14830 11398 14832 11450
rect 15012 11398 15014 11450
rect 14768 11396 14774 11398
rect 14830 11396 14854 11398
rect 14910 11396 14934 11398
rect 14990 11396 15014 11398
rect 15070 11396 15076 11398
rect 14768 11387 15076 11396
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 13912 10736 13964 10742
rect 13818 10704 13874 10713
rect 13912 10678 13964 10684
rect 13818 10639 13820 10648
rect 13872 10639 13874 10648
rect 13820 10610 13872 10616
rect 14108 10266 14136 10746
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14476 10169 14504 10406
rect 14462 10160 14518 10169
rect 14462 10095 14518 10104
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14292 9382 14320 9998
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14660 8430 14688 10610
rect 14768 10364 15076 10373
rect 14768 10362 14774 10364
rect 14830 10362 14854 10364
rect 14910 10362 14934 10364
rect 14990 10362 15014 10364
rect 15070 10362 15076 10364
rect 14830 10310 14832 10362
rect 15012 10310 15014 10362
rect 14768 10308 14774 10310
rect 14830 10308 14854 10310
rect 14910 10308 14934 10310
rect 14990 10308 15014 10310
rect 15070 10308 15076 10310
rect 14768 10299 15076 10308
rect 14768 9276 15076 9285
rect 14768 9274 14774 9276
rect 14830 9274 14854 9276
rect 14910 9274 14934 9276
rect 14990 9274 15014 9276
rect 15070 9274 15076 9276
rect 14830 9222 14832 9274
rect 15012 9222 15014 9274
rect 14768 9220 14774 9222
rect 14830 9220 14854 9222
rect 14910 9220 14934 9222
rect 14990 9220 15014 9222
rect 15070 9220 15076 9222
rect 14768 9211 15076 9220
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14768 8188 15076 8197
rect 14768 8186 14774 8188
rect 14830 8186 14854 8188
rect 14910 8186 14934 8188
rect 14990 8186 15014 8188
rect 15070 8186 15076 8188
rect 14830 8134 14832 8186
rect 15012 8134 15014 8186
rect 14768 8132 14774 8134
rect 14830 8132 14854 8134
rect 14910 8132 14934 8134
rect 14990 8132 15014 8134
rect 15070 8132 15076 8134
rect 14768 8123 15076 8132
rect 13176 7958 13228 7964
rect 13542 7984 13598 7993
rect 13542 7919 13598 7928
rect 12794 7644 13102 7653
rect 12794 7642 12800 7644
rect 12856 7642 12880 7644
rect 12936 7642 12960 7644
rect 13016 7642 13040 7644
rect 13096 7642 13102 7644
rect 12856 7590 12858 7642
rect 13038 7590 13040 7642
rect 12794 7588 12800 7590
rect 12856 7588 12880 7590
rect 12936 7588 12960 7590
rect 13016 7588 13040 7590
rect 13096 7588 13102 7590
rect 12794 7579 13102 7588
rect 14768 7100 15076 7109
rect 14768 7098 14774 7100
rect 14830 7098 14854 7100
rect 14910 7098 14934 7100
rect 14990 7098 15014 7100
rect 15070 7098 15076 7100
rect 14830 7046 14832 7098
rect 15012 7046 15014 7098
rect 14768 7044 14774 7046
rect 14830 7044 14854 7046
rect 14910 7044 14934 7046
rect 14990 7044 15014 7046
rect 15070 7044 15076 7046
rect 14768 7035 15076 7044
rect 12714 6760 12770 6769
rect 12714 6695 12770 6704
rect 12794 6556 13102 6565
rect 12794 6554 12800 6556
rect 12856 6554 12880 6556
rect 12936 6554 12960 6556
rect 13016 6554 13040 6556
rect 13096 6554 13102 6556
rect 12856 6502 12858 6554
rect 13038 6502 13040 6554
rect 12794 6500 12800 6502
rect 12856 6500 12880 6502
rect 12936 6500 12960 6502
rect 13016 6500 13040 6502
rect 13096 6500 13102 6502
rect 12794 6491 13102 6500
rect 14768 6012 15076 6021
rect 14768 6010 14774 6012
rect 14830 6010 14854 6012
rect 14910 6010 14934 6012
rect 14990 6010 15014 6012
rect 15070 6010 15076 6012
rect 14830 5958 14832 6010
rect 15012 5958 15014 6010
rect 14768 5956 14774 5958
rect 14830 5956 14854 5958
rect 14910 5956 14934 5958
rect 14990 5956 15014 5958
rect 15070 5956 15076 5958
rect 14768 5947 15076 5956
rect 12794 5468 13102 5477
rect 12794 5466 12800 5468
rect 12856 5466 12880 5468
rect 12936 5466 12960 5468
rect 13016 5466 13040 5468
rect 13096 5466 13102 5468
rect 12856 5414 12858 5466
rect 13038 5414 13040 5466
rect 12794 5412 12800 5414
rect 12856 5412 12880 5414
rect 12936 5412 12960 5414
rect 13016 5412 13040 5414
rect 13096 5412 13102 5414
rect 12794 5403 13102 5412
rect 14768 4924 15076 4933
rect 14768 4922 14774 4924
rect 14830 4922 14854 4924
rect 14910 4922 14934 4924
rect 14990 4922 15014 4924
rect 15070 4922 15076 4924
rect 14830 4870 14832 4922
rect 15012 4870 15014 4922
rect 14768 4868 14774 4870
rect 14830 4868 14854 4870
rect 14910 4868 14934 4870
rect 14990 4868 15014 4870
rect 15070 4868 15076 4870
rect 14768 4859 15076 4868
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12794 4380 13102 4389
rect 12794 4378 12800 4380
rect 12856 4378 12880 4380
rect 12936 4378 12960 4380
rect 13016 4378 13040 4380
rect 13096 4378 13102 4380
rect 12856 4326 12858 4378
rect 13038 4326 13040 4378
rect 12794 4324 12800 4326
rect 12856 4324 12880 4326
rect 12936 4324 12960 4326
rect 13016 4324 13040 4326
rect 13096 4324 13102 4326
rect 12794 4315 13102 4324
rect 14768 3836 15076 3845
rect 14768 3834 14774 3836
rect 14830 3834 14854 3836
rect 14910 3834 14934 3836
rect 14990 3834 15014 3836
rect 15070 3834 15076 3836
rect 14830 3782 14832 3834
rect 15012 3782 15014 3834
rect 14768 3780 14774 3782
rect 14830 3780 14854 3782
rect 14910 3780 14934 3782
rect 14990 3780 15014 3782
rect 15070 3780 15076 3782
rect 14768 3771 15076 3780
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 12794 3292 13102 3301
rect 12794 3290 12800 3292
rect 12856 3290 12880 3292
rect 12936 3290 12960 3292
rect 13016 3290 13040 3292
rect 13096 3290 13102 3292
rect 12856 3238 12858 3290
rect 13038 3238 13040 3290
rect 12794 3236 12800 3238
rect 12856 3236 12880 3238
rect 12936 3236 12960 3238
rect 13016 3236 13040 3238
rect 13096 3236 13102 3238
rect 12794 3227 13102 3236
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 6872 2748 7180 2757
rect 6872 2746 6878 2748
rect 6934 2746 6958 2748
rect 7014 2746 7038 2748
rect 7094 2746 7118 2748
rect 7174 2746 7180 2748
rect 6934 2694 6936 2746
rect 7116 2694 7118 2746
rect 6872 2692 6878 2694
rect 6934 2692 6958 2694
rect 7014 2692 7038 2694
rect 7094 2692 7118 2694
rect 7174 2692 7180 2694
rect 6872 2683 7180 2692
rect 10820 2748 11128 2757
rect 10820 2746 10826 2748
rect 10882 2746 10906 2748
rect 10962 2746 10986 2748
rect 11042 2746 11066 2748
rect 11122 2746 11128 2748
rect 10882 2694 10884 2746
rect 11064 2694 11066 2746
rect 10820 2692 10826 2694
rect 10882 2692 10906 2694
rect 10962 2692 10986 2694
rect 11042 2692 11066 2694
rect 11122 2692 11128 2694
rect 10820 2683 11128 2692
rect 14768 2748 15076 2757
rect 14768 2746 14774 2748
rect 14830 2746 14854 2748
rect 14910 2746 14934 2748
rect 14990 2746 15014 2748
rect 15070 2746 15076 2748
rect 14830 2694 14832 2746
rect 15012 2694 15014 2746
rect 14768 2692 14774 2694
rect 14830 2692 14854 2694
rect 14910 2692 14934 2694
rect 14990 2692 15014 2694
rect 15070 2692 15076 2694
rect 14768 2683 15076 2692
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 4898 2204 5206 2213
rect 4898 2202 4904 2204
rect 4960 2202 4984 2204
rect 5040 2202 5064 2204
rect 5120 2202 5144 2204
rect 5200 2202 5206 2204
rect 4960 2150 4962 2202
rect 5142 2150 5144 2202
rect 4898 2148 4904 2150
rect 4960 2148 4984 2150
rect 5040 2148 5064 2150
rect 5120 2148 5144 2150
rect 5200 2148 5206 2150
rect 4898 2139 5206 2148
rect 8846 2204 9154 2213
rect 8846 2202 8852 2204
rect 8908 2202 8932 2204
rect 8988 2202 9012 2204
rect 9068 2202 9092 2204
rect 9148 2202 9154 2204
rect 8908 2150 8910 2202
rect 9090 2150 9092 2202
rect 8846 2148 8852 2150
rect 8908 2148 8932 2150
rect 8988 2148 9012 2150
rect 9068 2148 9092 2150
rect 9148 2148 9154 2150
rect 8846 2139 9154 2148
rect 12794 2204 13102 2213
rect 12794 2202 12800 2204
rect 12856 2202 12880 2204
rect 12936 2202 12960 2204
rect 13016 2202 13040 2204
rect 13096 2202 13102 2204
rect 12856 2150 12858 2202
rect 13038 2150 13040 2202
rect 12794 2148 12800 2150
rect 12856 2148 12880 2150
rect 12936 2148 12960 2150
rect 13016 2148 13040 2150
rect 13096 2148 13102 2150
rect 12794 2139 13102 2148
rect 3608 2100 3660 2106
rect 3608 2042 3660 2048
rect 3424 2032 3476 2038
rect 3424 1974 3476 1980
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 2924 1660 3232 1669
rect 2924 1658 2930 1660
rect 2986 1658 3010 1660
rect 3066 1658 3090 1660
rect 3146 1658 3170 1660
rect 3226 1658 3232 1660
rect 2986 1606 2988 1658
rect 3168 1606 3170 1658
rect 2924 1604 2930 1606
rect 2986 1604 3010 1606
rect 3066 1604 3090 1606
rect 3146 1604 3170 1606
rect 3226 1604 3232 1606
rect 2924 1595 3232 1604
rect 6872 1660 7180 1669
rect 6872 1658 6878 1660
rect 6934 1658 6958 1660
rect 7014 1658 7038 1660
rect 7094 1658 7118 1660
rect 7174 1658 7180 1660
rect 6934 1606 6936 1658
rect 7116 1606 7118 1658
rect 6872 1604 6878 1606
rect 6934 1604 6958 1606
rect 7014 1604 7038 1606
rect 7094 1604 7118 1606
rect 7174 1604 7180 1606
rect 6872 1595 7180 1604
rect 10820 1660 11128 1669
rect 10820 1658 10826 1660
rect 10882 1658 10906 1660
rect 10962 1658 10986 1660
rect 11042 1658 11066 1660
rect 11122 1658 11128 1660
rect 10882 1606 10884 1658
rect 11064 1606 11066 1658
rect 10820 1604 10826 1606
rect 10882 1604 10906 1606
rect 10962 1604 10986 1606
rect 11042 1604 11066 1606
rect 11122 1604 11128 1606
rect 10820 1595 11128 1604
rect 14768 1660 15076 1669
rect 14768 1658 14774 1660
rect 14830 1658 14854 1660
rect 14910 1658 14934 1660
rect 14990 1658 15014 1660
rect 15070 1658 15076 1660
rect 14830 1606 14832 1658
rect 15012 1606 15014 1658
rect 14768 1604 14774 1606
rect 14830 1604 14854 1606
rect 14910 1604 14934 1606
rect 14990 1604 15014 1606
rect 15070 1604 15076 1606
rect 14768 1595 15076 1604
rect 1492 1216 1544 1222
rect 1492 1158 1544 1164
rect 4898 1116 5206 1125
rect 4898 1114 4904 1116
rect 4960 1114 4984 1116
rect 5040 1114 5064 1116
rect 5120 1114 5144 1116
rect 5200 1114 5206 1116
rect 4960 1062 4962 1114
rect 5142 1062 5144 1114
rect 4898 1060 4904 1062
rect 4960 1060 4984 1062
rect 5040 1060 5064 1062
rect 5120 1060 5144 1062
rect 5200 1060 5206 1062
rect 4898 1051 5206 1060
rect 8846 1116 9154 1125
rect 8846 1114 8852 1116
rect 8908 1114 8932 1116
rect 8988 1114 9012 1116
rect 9068 1114 9092 1116
rect 9148 1114 9154 1116
rect 8908 1062 8910 1114
rect 9090 1062 9092 1114
rect 8846 1060 8852 1062
rect 8908 1060 8932 1062
rect 8988 1060 9012 1062
rect 9068 1060 9092 1062
rect 9148 1060 9154 1062
rect 8846 1051 9154 1060
rect 12794 1116 13102 1125
rect 12794 1114 12800 1116
rect 12856 1114 12880 1116
rect 12936 1114 12960 1116
rect 13016 1114 13040 1116
rect 13096 1114 13102 1116
rect 12856 1062 12858 1114
rect 13038 1062 13040 1114
rect 12794 1060 12800 1062
rect 12856 1060 12880 1062
rect 12936 1060 12960 1062
rect 13016 1060 13040 1062
rect 13096 1060 13102 1062
rect 12794 1051 13102 1060
rect 1398 776 1454 785
rect 1398 711 1454 720
<< via2 >>
rect 2778 23160 2834 23216
rect 1490 21664 1546 21720
rect 4904 22874 4960 22876
rect 4984 22874 5040 22876
rect 5064 22874 5120 22876
rect 5144 22874 5200 22876
rect 4904 22822 4950 22874
rect 4950 22822 4960 22874
rect 4984 22822 5014 22874
rect 5014 22822 5026 22874
rect 5026 22822 5040 22874
rect 5064 22822 5078 22874
rect 5078 22822 5090 22874
rect 5090 22822 5120 22874
rect 5144 22822 5154 22874
rect 5154 22822 5200 22874
rect 4904 22820 4960 22822
rect 4984 22820 5040 22822
rect 5064 22820 5120 22822
rect 5144 22820 5200 22822
rect 8852 22874 8908 22876
rect 8932 22874 8988 22876
rect 9012 22874 9068 22876
rect 9092 22874 9148 22876
rect 8852 22822 8898 22874
rect 8898 22822 8908 22874
rect 8932 22822 8962 22874
rect 8962 22822 8974 22874
rect 8974 22822 8988 22874
rect 9012 22822 9026 22874
rect 9026 22822 9038 22874
rect 9038 22822 9068 22874
rect 9092 22822 9102 22874
rect 9102 22822 9148 22874
rect 8852 22820 8908 22822
rect 8932 22820 8988 22822
rect 9012 22820 9068 22822
rect 9092 22820 9148 22822
rect 12800 22874 12856 22876
rect 12880 22874 12936 22876
rect 12960 22874 13016 22876
rect 13040 22874 13096 22876
rect 12800 22822 12846 22874
rect 12846 22822 12856 22874
rect 12880 22822 12910 22874
rect 12910 22822 12922 22874
rect 12922 22822 12936 22874
rect 12960 22822 12974 22874
rect 12974 22822 12986 22874
rect 12986 22822 13016 22874
rect 13040 22822 13050 22874
rect 13050 22822 13096 22874
rect 12800 22820 12856 22822
rect 12880 22820 12936 22822
rect 12960 22820 13016 22822
rect 13040 22820 13096 22822
rect 2930 22330 2986 22332
rect 3010 22330 3066 22332
rect 3090 22330 3146 22332
rect 3170 22330 3226 22332
rect 2930 22278 2976 22330
rect 2976 22278 2986 22330
rect 3010 22278 3040 22330
rect 3040 22278 3052 22330
rect 3052 22278 3066 22330
rect 3090 22278 3104 22330
rect 3104 22278 3116 22330
rect 3116 22278 3146 22330
rect 3170 22278 3180 22330
rect 3180 22278 3226 22330
rect 2930 22276 2986 22278
rect 3010 22276 3066 22278
rect 3090 22276 3146 22278
rect 3170 22276 3226 22278
rect 6878 22330 6934 22332
rect 6958 22330 7014 22332
rect 7038 22330 7094 22332
rect 7118 22330 7174 22332
rect 6878 22278 6924 22330
rect 6924 22278 6934 22330
rect 6958 22278 6988 22330
rect 6988 22278 7000 22330
rect 7000 22278 7014 22330
rect 7038 22278 7052 22330
rect 7052 22278 7064 22330
rect 7064 22278 7094 22330
rect 7118 22278 7128 22330
rect 7128 22278 7174 22330
rect 6878 22276 6934 22278
rect 6958 22276 7014 22278
rect 7038 22276 7094 22278
rect 7118 22276 7174 22278
rect 10826 22330 10882 22332
rect 10906 22330 10962 22332
rect 10986 22330 11042 22332
rect 11066 22330 11122 22332
rect 10826 22278 10872 22330
rect 10872 22278 10882 22330
rect 10906 22278 10936 22330
rect 10936 22278 10948 22330
rect 10948 22278 10962 22330
rect 10986 22278 11000 22330
rect 11000 22278 11012 22330
rect 11012 22278 11042 22330
rect 11066 22278 11076 22330
rect 11076 22278 11122 22330
rect 10826 22276 10882 22278
rect 10906 22276 10962 22278
rect 10986 22276 11042 22278
rect 11066 22276 11122 22278
rect 14774 22330 14830 22332
rect 14854 22330 14910 22332
rect 14934 22330 14990 22332
rect 15014 22330 15070 22332
rect 14774 22278 14820 22330
rect 14820 22278 14830 22330
rect 14854 22278 14884 22330
rect 14884 22278 14896 22330
rect 14896 22278 14910 22330
rect 14934 22278 14948 22330
rect 14948 22278 14960 22330
rect 14960 22278 14990 22330
rect 15014 22278 15024 22330
rect 15024 22278 15070 22330
rect 14774 22276 14830 22278
rect 14854 22276 14910 22278
rect 14934 22276 14990 22278
rect 15014 22276 15070 22278
rect 4904 21786 4960 21788
rect 4984 21786 5040 21788
rect 5064 21786 5120 21788
rect 5144 21786 5200 21788
rect 4904 21734 4950 21786
rect 4950 21734 4960 21786
rect 4984 21734 5014 21786
rect 5014 21734 5026 21786
rect 5026 21734 5040 21786
rect 5064 21734 5078 21786
rect 5078 21734 5090 21786
rect 5090 21734 5120 21786
rect 5144 21734 5154 21786
rect 5154 21734 5200 21786
rect 4904 21732 4960 21734
rect 4984 21732 5040 21734
rect 5064 21732 5120 21734
rect 5144 21732 5200 21734
rect 8852 21786 8908 21788
rect 8932 21786 8988 21788
rect 9012 21786 9068 21788
rect 9092 21786 9148 21788
rect 8852 21734 8898 21786
rect 8898 21734 8908 21786
rect 8932 21734 8962 21786
rect 8962 21734 8974 21786
rect 8974 21734 8988 21786
rect 9012 21734 9026 21786
rect 9026 21734 9038 21786
rect 9038 21734 9068 21786
rect 9092 21734 9102 21786
rect 9102 21734 9148 21786
rect 8852 21732 8908 21734
rect 8932 21732 8988 21734
rect 9012 21732 9068 21734
rect 9092 21732 9148 21734
rect 12800 21786 12856 21788
rect 12880 21786 12936 21788
rect 12960 21786 13016 21788
rect 13040 21786 13096 21788
rect 12800 21734 12846 21786
rect 12846 21734 12856 21786
rect 12880 21734 12910 21786
rect 12910 21734 12922 21786
rect 12922 21734 12936 21786
rect 12960 21734 12974 21786
rect 12974 21734 12986 21786
rect 12986 21734 13016 21786
rect 13040 21734 13050 21786
rect 13050 21734 13096 21786
rect 12800 21732 12856 21734
rect 12880 21732 12936 21734
rect 12960 21732 13016 21734
rect 13040 21732 13096 21734
rect 2930 21242 2986 21244
rect 3010 21242 3066 21244
rect 3090 21242 3146 21244
rect 3170 21242 3226 21244
rect 2930 21190 2976 21242
rect 2976 21190 2986 21242
rect 3010 21190 3040 21242
rect 3040 21190 3052 21242
rect 3052 21190 3066 21242
rect 3090 21190 3104 21242
rect 3104 21190 3116 21242
rect 3116 21190 3146 21242
rect 3170 21190 3180 21242
rect 3180 21190 3226 21242
rect 2930 21188 2986 21190
rect 3010 21188 3066 21190
rect 3090 21188 3146 21190
rect 3170 21188 3226 21190
rect 6878 21242 6934 21244
rect 6958 21242 7014 21244
rect 7038 21242 7094 21244
rect 7118 21242 7174 21244
rect 6878 21190 6924 21242
rect 6924 21190 6934 21242
rect 6958 21190 6988 21242
rect 6988 21190 7000 21242
rect 7000 21190 7014 21242
rect 7038 21190 7052 21242
rect 7052 21190 7064 21242
rect 7064 21190 7094 21242
rect 7118 21190 7128 21242
rect 7128 21190 7174 21242
rect 6878 21188 6934 21190
rect 6958 21188 7014 21190
rect 7038 21188 7094 21190
rect 7118 21188 7174 21190
rect 10826 21242 10882 21244
rect 10906 21242 10962 21244
rect 10986 21242 11042 21244
rect 11066 21242 11122 21244
rect 10826 21190 10872 21242
rect 10872 21190 10882 21242
rect 10906 21190 10936 21242
rect 10936 21190 10948 21242
rect 10948 21190 10962 21242
rect 10986 21190 11000 21242
rect 11000 21190 11012 21242
rect 11012 21190 11042 21242
rect 11066 21190 11076 21242
rect 11076 21190 11122 21242
rect 10826 21188 10882 21190
rect 10906 21188 10962 21190
rect 10986 21188 11042 21190
rect 11066 21188 11122 21190
rect 14774 21242 14830 21244
rect 14854 21242 14910 21244
rect 14934 21242 14990 21244
rect 15014 21242 15070 21244
rect 14774 21190 14820 21242
rect 14820 21190 14830 21242
rect 14854 21190 14884 21242
rect 14884 21190 14896 21242
rect 14896 21190 14910 21242
rect 14934 21190 14948 21242
rect 14948 21190 14960 21242
rect 14960 21190 14990 21242
rect 15014 21190 15024 21242
rect 15024 21190 15070 21242
rect 14774 21188 14830 21190
rect 14854 21188 14910 21190
rect 14934 21188 14990 21190
rect 15014 21188 15070 21190
rect 4904 20698 4960 20700
rect 4984 20698 5040 20700
rect 5064 20698 5120 20700
rect 5144 20698 5200 20700
rect 4904 20646 4950 20698
rect 4950 20646 4960 20698
rect 4984 20646 5014 20698
rect 5014 20646 5026 20698
rect 5026 20646 5040 20698
rect 5064 20646 5078 20698
rect 5078 20646 5090 20698
rect 5090 20646 5120 20698
rect 5144 20646 5154 20698
rect 5154 20646 5200 20698
rect 4904 20644 4960 20646
rect 4984 20644 5040 20646
rect 5064 20644 5120 20646
rect 5144 20644 5200 20646
rect 8852 20698 8908 20700
rect 8932 20698 8988 20700
rect 9012 20698 9068 20700
rect 9092 20698 9148 20700
rect 8852 20646 8898 20698
rect 8898 20646 8908 20698
rect 8932 20646 8962 20698
rect 8962 20646 8974 20698
rect 8974 20646 8988 20698
rect 9012 20646 9026 20698
rect 9026 20646 9038 20698
rect 9038 20646 9068 20698
rect 9092 20646 9102 20698
rect 9102 20646 9148 20698
rect 8852 20644 8908 20646
rect 8932 20644 8988 20646
rect 9012 20644 9068 20646
rect 9092 20644 9148 20646
rect 12800 20698 12856 20700
rect 12880 20698 12936 20700
rect 12960 20698 13016 20700
rect 13040 20698 13096 20700
rect 12800 20646 12846 20698
rect 12846 20646 12856 20698
rect 12880 20646 12910 20698
rect 12910 20646 12922 20698
rect 12922 20646 12936 20698
rect 12960 20646 12974 20698
rect 12974 20646 12986 20698
rect 12986 20646 13016 20698
rect 13040 20646 13050 20698
rect 13050 20646 13096 20698
rect 12800 20644 12856 20646
rect 12880 20644 12936 20646
rect 12960 20644 13016 20646
rect 13040 20644 13096 20646
rect 2930 20154 2986 20156
rect 3010 20154 3066 20156
rect 3090 20154 3146 20156
rect 3170 20154 3226 20156
rect 2930 20102 2976 20154
rect 2976 20102 2986 20154
rect 3010 20102 3040 20154
rect 3040 20102 3052 20154
rect 3052 20102 3066 20154
rect 3090 20102 3104 20154
rect 3104 20102 3116 20154
rect 3116 20102 3146 20154
rect 3170 20102 3180 20154
rect 3180 20102 3226 20154
rect 2930 20100 2986 20102
rect 3010 20100 3066 20102
rect 3090 20100 3146 20102
rect 3170 20100 3226 20102
rect 6878 20154 6934 20156
rect 6958 20154 7014 20156
rect 7038 20154 7094 20156
rect 7118 20154 7174 20156
rect 6878 20102 6924 20154
rect 6924 20102 6934 20154
rect 6958 20102 6988 20154
rect 6988 20102 7000 20154
rect 7000 20102 7014 20154
rect 7038 20102 7052 20154
rect 7052 20102 7064 20154
rect 7064 20102 7094 20154
rect 7118 20102 7128 20154
rect 7128 20102 7174 20154
rect 6878 20100 6934 20102
rect 6958 20100 7014 20102
rect 7038 20100 7094 20102
rect 7118 20100 7174 20102
rect 10826 20154 10882 20156
rect 10906 20154 10962 20156
rect 10986 20154 11042 20156
rect 11066 20154 11122 20156
rect 10826 20102 10872 20154
rect 10872 20102 10882 20154
rect 10906 20102 10936 20154
rect 10936 20102 10948 20154
rect 10948 20102 10962 20154
rect 10986 20102 11000 20154
rect 11000 20102 11012 20154
rect 11012 20102 11042 20154
rect 11066 20102 11076 20154
rect 11076 20102 11122 20154
rect 10826 20100 10882 20102
rect 10906 20100 10962 20102
rect 10986 20100 11042 20102
rect 11066 20100 11122 20102
rect 14774 20154 14830 20156
rect 14854 20154 14910 20156
rect 14934 20154 14990 20156
rect 15014 20154 15070 20156
rect 14774 20102 14820 20154
rect 14820 20102 14830 20154
rect 14854 20102 14884 20154
rect 14884 20102 14896 20154
rect 14896 20102 14910 20154
rect 14934 20102 14948 20154
rect 14948 20102 14960 20154
rect 14960 20102 14990 20154
rect 15014 20102 15024 20154
rect 15024 20102 15070 20154
rect 14774 20100 14830 20102
rect 14854 20100 14910 20102
rect 14934 20100 14990 20102
rect 15014 20100 15070 20102
rect 3330 19896 3386 19952
rect 2930 19066 2986 19068
rect 3010 19066 3066 19068
rect 3090 19066 3146 19068
rect 3170 19066 3226 19068
rect 2930 19014 2976 19066
rect 2976 19014 2986 19066
rect 3010 19014 3040 19066
rect 3040 19014 3052 19066
rect 3052 19014 3066 19066
rect 3090 19014 3104 19066
rect 3104 19014 3116 19066
rect 3116 19014 3146 19066
rect 3170 19014 3180 19066
rect 3180 19014 3226 19066
rect 2930 19012 2986 19014
rect 3010 19012 3066 19014
rect 3090 19012 3146 19014
rect 3170 19012 3226 19014
rect 2778 18672 2834 18728
rect 1490 17176 1546 17232
rect 2042 14864 2098 14920
rect 2930 17978 2986 17980
rect 3010 17978 3066 17980
rect 3090 17978 3146 17980
rect 3170 17978 3226 17980
rect 2930 17926 2976 17978
rect 2976 17926 2986 17978
rect 3010 17926 3040 17978
rect 3040 17926 3052 17978
rect 3052 17926 3066 17978
rect 3090 17926 3104 17978
rect 3104 17926 3116 17978
rect 3116 17926 3146 17978
rect 3170 17926 3180 17978
rect 3180 17926 3226 17978
rect 2930 17924 2986 17926
rect 3010 17924 3066 17926
rect 3090 17924 3146 17926
rect 3170 17924 3226 17926
rect 4904 19610 4960 19612
rect 4984 19610 5040 19612
rect 5064 19610 5120 19612
rect 5144 19610 5200 19612
rect 4904 19558 4950 19610
rect 4950 19558 4960 19610
rect 4984 19558 5014 19610
rect 5014 19558 5026 19610
rect 5026 19558 5040 19610
rect 5064 19558 5078 19610
rect 5078 19558 5090 19610
rect 5090 19558 5120 19610
rect 5144 19558 5154 19610
rect 5154 19558 5200 19610
rect 4904 19556 4960 19558
rect 4984 19556 5040 19558
rect 5064 19556 5120 19558
rect 5144 19556 5200 19558
rect 8852 19610 8908 19612
rect 8932 19610 8988 19612
rect 9012 19610 9068 19612
rect 9092 19610 9148 19612
rect 8852 19558 8898 19610
rect 8898 19558 8908 19610
rect 8932 19558 8962 19610
rect 8962 19558 8974 19610
rect 8974 19558 8988 19610
rect 9012 19558 9026 19610
rect 9026 19558 9038 19610
rect 9038 19558 9068 19610
rect 9092 19558 9102 19610
rect 9102 19558 9148 19610
rect 8852 19556 8908 19558
rect 8932 19556 8988 19558
rect 9012 19556 9068 19558
rect 9092 19556 9148 19558
rect 12800 19610 12856 19612
rect 12880 19610 12936 19612
rect 12960 19610 13016 19612
rect 13040 19610 13096 19612
rect 12800 19558 12846 19610
rect 12846 19558 12856 19610
rect 12880 19558 12910 19610
rect 12910 19558 12922 19610
rect 12922 19558 12936 19610
rect 12960 19558 12974 19610
rect 12974 19558 12986 19610
rect 12986 19558 13016 19610
rect 13040 19558 13050 19610
rect 13050 19558 13096 19610
rect 12800 19556 12856 19558
rect 12880 19556 12936 19558
rect 12960 19556 13016 19558
rect 13040 19556 13096 19558
rect 6878 19066 6934 19068
rect 6958 19066 7014 19068
rect 7038 19066 7094 19068
rect 7118 19066 7174 19068
rect 6878 19014 6924 19066
rect 6924 19014 6934 19066
rect 6958 19014 6988 19066
rect 6988 19014 7000 19066
rect 7000 19014 7014 19066
rect 7038 19014 7052 19066
rect 7052 19014 7064 19066
rect 7064 19014 7094 19066
rect 7118 19014 7128 19066
rect 7128 19014 7174 19066
rect 6878 19012 6934 19014
rect 6958 19012 7014 19014
rect 7038 19012 7094 19014
rect 7118 19012 7174 19014
rect 10826 19066 10882 19068
rect 10906 19066 10962 19068
rect 10986 19066 11042 19068
rect 11066 19066 11122 19068
rect 10826 19014 10872 19066
rect 10872 19014 10882 19066
rect 10906 19014 10936 19066
rect 10936 19014 10948 19066
rect 10948 19014 10962 19066
rect 10986 19014 11000 19066
rect 11000 19014 11012 19066
rect 11012 19014 11042 19066
rect 11066 19014 11076 19066
rect 11076 19014 11122 19066
rect 10826 19012 10882 19014
rect 10906 19012 10962 19014
rect 10986 19012 11042 19014
rect 11066 19012 11122 19014
rect 14774 19066 14830 19068
rect 14854 19066 14910 19068
rect 14934 19066 14990 19068
rect 15014 19066 15070 19068
rect 14774 19014 14820 19066
rect 14820 19014 14830 19066
rect 14854 19014 14884 19066
rect 14884 19014 14896 19066
rect 14896 19014 14910 19066
rect 14934 19014 14948 19066
rect 14948 19014 14960 19066
rect 14960 19014 14990 19066
rect 15014 19014 15024 19066
rect 15024 19014 15070 19066
rect 14774 19012 14830 19014
rect 14854 19012 14910 19014
rect 14934 19012 14990 19014
rect 15014 19012 15070 19014
rect 2930 16890 2986 16892
rect 3010 16890 3066 16892
rect 3090 16890 3146 16892
rect 3170 16890 3226 16892
rect 2930 16838 2976 16890
rect 2976 16838 2986 16890
rect 3010 16838 3040 16890
rect 3040 16838 3052 16890
rect 3052 16838 3066 16890
rect 3090 16838 3104 16890
rect 3104 16838 3116 16890
rect 3116 16838 3146 16890
rect 3170 16838 3180 16890
rect 3180 16838 3226 16890
rect 2930 16836 2986 16838
rect 3010 16836 3066 16838
rect 3090 16836 3146 16838
rect 3170 16836 3226 16838
rect 2930 15802 2986 15804
rect 3010 15802 3066 15804
rect 3090 15802 3146 15804
rect 3170 15802 3226 15804
rect 2930 15750 2976 15802
rect 2976 15750 2986 15802
rect 3010 15750 3040 15802
rect 3040 15750 3052 15802
rect 3052 15750 3066 15802
rect 3090 15750 3104 15802
rect 3104 15750 3116 15802
rect 3116 15750 3146 15802
rect 3170 15750 3180 15802
rect 3180 15750 3226 15802
rect 2930 15748 2986 15750
rect 3010 15748 3066 15750
rect 3090 15748 3146 15750
rect 3170 15748 3226 15750
rect 2778 15680 2834 15736
rect 2930 14714 2986 14716
rect 3010 14714 3066 14716
rect 3090 14714 3146 14716
rect 3170 14714 3226 14716
rect 2930 14662 2976 14714
rect 2976 14662 2986 14714
rect 3010 14662 3040 14714
rect 3040 14662 3052 14714
rect 3052 14662 3066 14714
rect 3090 14662 3104 14714
rect 3104 14662 3116 14714
rect 3116 14662 3146 14714
rect 3170 14662 3180 14714
rect 3180 14662 3226 14714
rect 2930 14660 2986 14662
rect 3010 14660 3066 14662
rect 3090 14660 3146 14662
rect 3170 14660 3226 14662
rect 3422 15000 3478 15056
rect 3330 14184 3386 14240
rect 2930 13626 2986 13628
rect 3010 13626 3066 13628
rect 3090 13626 3146 13628
rect 3170 13626 3226 13628
rect 2930 13574 2976 13626
rect 2976 13574 2986 13626
rect 3010 13574 3040 13626
rect 3040 13574 3052 13626
rect 3052 13574 3066 13626
rect 3090 13574 3104 13626
rect 3104 13574 3116 13626
rect 3116 13574 3146 13626
rect 3170 13574 3180 13626
rect 3180 13574 3226 13626
rect 2930 13572 2986 13574
rect 3010 13572 3066 13574
rect 3090 13572 3146 13574
rect 3170 13572 3226 13574
rect 2686 13368 2742 13424
rect 2778 13232 2834 13288
rect 2962 12844 3018 12880
rect 2962 12824 2964 12844
rect 2964 12824 3016 12844
rect 3016 12824 3018 12844
rect 2930 12538 2986 12540
rect 3010 12538 3066 12540
rect 3090 12538 3146 12540
rect 3170 12538 3226 12540
rect 2930 12486 2976 12538
rect 2976 12486 2986 12538
rect 3010 12486 3040 12538
rect 3040 12486 3052 12538
rect 3052 12486 3066 12538
rect 3090 12486 3104 12538
rect 3104 12486 3116 12538
rect 3116 12486 3146 12538
rect 3170 12486 3180 12538
rect 3180 12486 3226 12538
rect 2930 12484 2986 12486
rect 3010 12484 3066 12486
rect 3090 12484 3146 12486
rect 3170 12484 3226 12486
rect 2502 12300 2558 12336
rect 2502 12280 2504 12300
rect 2504 12280 2556 12300
rect 2556 12280 2558 12300
rect 3514 12688 3570 12744
rect 3422 12552 3478 12608
rect 4342 15544 4398 15600
rect 4904 18522 4960 18524
rect 4984 18522 5040 18524
rect 5064 18522 5120 18524
rect 5144 18522 5200 18524
rect 4904 18470 4950 18522
rect 4950 18470 4960 18522
rect 4984 18470 5014 18522
rect 5014 18470 5026 18522
rect 5026 18470 5040 18522
rect 5064 18470 5078 18522
rect 5078 18470 5090 18522
rect 5090 18470 5120 18522
rect 5144 18470 5154 18522
rect 5154 18470 5200 18522
rect 4904 18468 4960 18470
rect 4984 18468 5040 18470
rect 5064 18468 5120 18470
rect 5144 18468 5200 18470
rect 8852 18522 8908 18524
rect 8932 18522 8988 18524
rect 9012 18522 9068 18524
rect 9092 18522 9148 18524
rect 8852 18470 8898 18522
rect 8898 18470 8908 18522
rect 8932 18470 8962 18522
rect 8962 18470 8974 18522
rect 8974 18470 8988 18522
rect 9012 18470 9026 18522
rect 9026 18470 9038 18522
rect 9038 18470 9068 18522
rect 9092 18470 9102 18522
rect 9102 18470 9148 18522
rect 8852 18468 8908 18470
rect 8932 18468 8988 18470
rect 9012 18468 9068 18470
rect 9092 18468 9148 18470
rect 12800 18522 12856 18524
rect 12880 18522 12936 18524
rect 12960 18522 13016 18524
rect 13040 18522 13096 18524
rect 12800 18470 12846 18522
rect 12846 18470 12856 18522
rect 12880 18470 12910 18522
rect 12910 18470 12922 18522
rect 12922 18470 12936 18522
rect 12960 18470 12974 18522
rect 12974 18470 12986 18522
rect 12986 18470 13016 18522
rect 13040 18470 13050 18522
rect 13050 18470 13096 18522
rect 12800 18468 12856 18470
rect 12880 18468 12936 18470
rect 12960 18468 13016 18470
rect 13040 18468 13096 18470
rect 6878 17978 6934 17980
rect 6958 17978 7014 17980
rect 7038 17978 7094 17980
rect 7118 17978 7174 17980
rect 6878 17926 6924 17978
rect 6924 17926 6934 17978
rect 6958 17926 6988 17978
rect 6988 17926 7000 17978
rect 7000 17926 7014 17978
rect 7038 17926 7052 17978
rect 7052 17926 7064 17978
rect 7064 17926 7094 17978
rect 7118 17926 7128 17978
rect 7128 17926 7174 17978
rect 6878 17924 6934 17926
rect 6958 17924 7014 17926
rect 7038 17924 7094 17926
rect 7118 17924 7174 17926
rect 10826 17978 10882 17980
rect 10906 17978 10962 17980
rect 10986 17978 11042 17980
rect 11066 17978 11122 17980
rect 10826 17926 10872 17978
rect 10872 17926 10882 17978
rect 10906 17926 10936 17978
rect 10936 17926 10948 17978
rect 10948 17926 10962 17978
rect 10986 17926 11000 17978
rect 11000 17926 11012 17978
rect 11012 17926 11042 17978
rect 11066 17926 11076 17978
rect 11076 17926 11122 17978
rect 10826 17924 10882 17926
rect 10906 17924 10962 17926
rect 10986 17924 11042 17926
rect 11066 17924 11122 17926
rect 14774 17978 14830 17980
rect 14854 17978 14910 17980
rect 14934 17978 14990 17980
rect 15014 17978 15070 17980
rect 14774 17926 14820 17978
rect 14820 17926 14830 17978
rect 14854 17926 14884 17978
rect 14884 17926 14896 17978
rect 14896 17926 14910 17978
rect 14934 17926 14948 17978
rect 14948 17926 14960 17978
rect 14960 17926 14990 17978
rect 15014 17926 15024 17978
rect 15024 17926 15070 17978
rect 14774 17924 14830 17926
rect 14854 17924 14910 17926
rect 14934 17924 14990 17926
rect 15014 17924 15070 17926
rect 4904 17434 4960 17436
rect 4984 17434 5040 17436
rect 5064 17434 5120 17436
rect 5144 17434 5200 17436
rect 4904 17382 4950 17434
rect 4950 17382 4960 17434
rect 4984 17382 5014 17434
rect 5014 17382 5026 17434
rect 5026 17382 5040 17434
rect 5064 17382 5078 17434
rect 5078 17382 5090 17434
rect 5090 17382 5120 17434
rect 5144 17382 5154 17434
rect 5154 17382 5200 17434
rect 4904 17380 4960 17382
rect 4984 17380 5040 17382
rect 5064 17380 5120 17382
rect 5144 17380 5200 17382
rect 8852 17434 8908 17436
rect 8932 17434 8988 17436
rect 9012 17434 9068 17436
rect 9092 17434 9148 17436
rect 8852 17382 8898 17434
rect 8898 17382 8908 17434
rect 8932 17382 8962 17434
rect 8962 17382 8974 17434
rect 8974 17382 8988 17434
rect 9012 17382 9026 17434
rect 9026 17382 9038 17434
rect 9038 17382 9068 17434
rect 9092 17382 9102 17434
rect 9102 17382 9148 17434
rect 8852 17380 8908 17382
rect 8932 17380 8988 17382
rect 9012 17380 9068 17382
rect 9092 17380 9148 17382
rect 12800 17434 12856 17436
rect 12880 17434 12936 17436
rect 12960 17434 13016 17436
rect 13040 17434 13096 17436
rect 12800 17382 12846 17434
rect 12846 17382 12856 17434
rect 12880 17382 12910 17434
rect 12910 17382 12922 17434
rect 12922 17382 12936 17434
rect 12960 17382 12974 17434
rect 12974 17382 12986 17434
rect 12986 17382 13016 17434
rect 13040 17382 13050 17434
rect 13050 17382 13096 17434
rect 12800 17380 12856 17382
rect 12880 17380 12936 17382
rect 12960 17380 13016 17382
rect 13040 17380 13096 17382
rect 4904 16346 4960 16348
rect 4984 16346 5040 16348
rect 5064 16346 5120 16348
rect 5144 16346 5200 16348
rect 4904 16294 4950 16346
rect 4950 16294 4960 16346
rect 4984 16294 5014 16346
rect 5014 16294 5026 16346
rect 5026 16294 5040 16346
rect 5064 16294 5078 16346
rect 5078 16294 5090 16346
rect 5090 16294 5120 16346
rect 5144 16294 5154 16346
rect 5154 16294 5200 16346
rect 4904 16292 4960 16294
rect 4984 16292 5040 16294
rect 5064 16292 5120 16294
rect 5144 16292 5200 16294
rect 3882 13504 3938 13560
rect 2930 11450 2986 11452
rect 3010 11450 3066 11452
rect 3090 11450 3146 11452
rect 3170 11450 3226 11452
rect 2930 11398 2976 11450
rect 2976 11398 2986 11450
rect 3010 11398 3040 11450
rect 3040 11398 3052 11450
rect 3052 11398 3066 11450
rect 3090 11398 3104 11450
rect 3104 11398 3116 11450
rect 3116 11398 3146 11450
rect 3170 11398 3180 11450
rect 3180 11398 3226 11450
rect 2930 11396 2986 11398
rect 3010 11396 3066 11398
rect 3090 11396 3146 11398
rect 3170 11396 3226 11398
rect 2778 10648 2834 10704
rect 1306 9424 1362 9480
rect 1490 9016 1546 9072
rect 2502 10512 2558 10568
rect 2930 10362 2986 10364
rect 3010 10362 3066 10364
rect 3090 10362 3146 10364
rect 3170 10362 3226 10364
rect 2930 10310 2976 10362
rect 2976 10310 2986 10362
rect 3010 10310 3040 10362
rect 3040 10310 3052 10362
rect 3052 10310 3066 10362
rect 3090 10310 3104 10362
rect 3104 10310 3116 10362
rect 3116 10310 3146 10362
rect 3170 10310 3180 10362
rect 3180 10310 3226 10362
rect 2930 10308 2986 10310
rect 3010 10308 3066 10310
rect 3090 10308 3146 10310
rect 3170 10308 3226 10310
rect 3422 10104 3478 10160
rect 1766 9988 1822 10024
rect 1766 9968 1768 9988
rect 1768 9968 1820 9988
rect 1820 9968 1822 9988
rect 2930 9274 2986 9276
rect 3010 9274 3066 9276
rect 3090 9274 3146 9276
rect 3170 9274 3226 9276
rect 2930 9222 2976 9274
rect 2976 9222 2986 9274
rect 3010 9222 3040 9274
rect 3040 9222 3052 9274
rect 3052 9222 3066 9274
rect 3090 9222 3104 9274
rect 3104 9222 3116 9274
rect 3116 9222 3146 9274
rect 3170 9222 3180 9274
rect 3180 9222 3226 9274
rect 2930 9220 2986 9222
rect 3010 9220 3066 9222
rect 3090 9220 3146 9222
rect 3170 9220 3226 9222
rect 2042 7792 2098 7848
rect 1398 6704 1454 6760
rect 1582 6160 1638 6216
rect 1490 4528 1546 4584
rect 1398 3712 1454 3768
rect 1306 3304 1362 3360
rect 1398 2216 1454 2272
rect 1858 7248 1914 7304
rect 1674 3984 1730 4040
rect 2686 8472 2742 8528
rect 2930 8186 2986 8188
rect 3010 8186 3066 8188
rect 3090 8186 3146 8188
rect 3170 8186 3226 8188
rect 2930 8134 2976 8186
rect 2976 8134 2986 8186
rect 3010 8134 3040 8186
rect 3040 8134 3052 8186
rect 3052 8134 3066 8186
rect 3090 8134 3104 8186
rect 3104 8134 3116 8186
rect 3116 8134 3146 8186
rect 3170 8134 3180 8186
rect 3180 8134 3226 8186
rect 2930 8132 2986 8134
rect 3010 8132 3066 8134
rect 3090 8132 3146 8134
rect 3170 8132 3226 8134
rect 2930 7098 2986 7100
rect 3010 7098 3066 7100
rect 3090 7098 3146 7100
rect 3170 7098 3226 7100
rect 2930 7046 2976 7098
rect 2976 7046 2986 7098
rect 3010 7046 3040 7098
rect 3040 7046 3052 7098
rect 3052 7046 3066 7098
rect 3090 7046 3104 7098
rect 3104 7046 3116 7098
rect 3116 7046 3146 7098
rect 3170 7046 3180 7098
rect 3180 7046 3226 7098
rect 2930 7044 2986 7046
rect 3010 7044 3066 7046
rect 3090 7044 3146 7046
rect 3170 7044 3226 7046
rect 2778 6296 2834 6352
rect 2930 6010 2986 6012
rect 3010 6010 3066 6012
rect 3090 6010 3146 6012
rect 3170 6010 3226 6012
rect 2930 5958 2976 6010
rect 2976 5958 2986 6010
rect 3010 5958 3040 6010
rect 3040 5958 3052 6010
rect 3052 5958 3066 6010
rect 3090 5958 3104 6010
rect 3104 5958 3116 6010
rect 3116 5958 3146 6010
rect 3170 5958 3180 6010
rect 3180 5958 3226 6010
rect 2930 5956 2986 5958
rect 3010 5956 3066 5958
rect 3090 5956 3146 5958
rect 3170 5956 3226 5958
rect 3054 5344 3110 5400
rect 2226 3052 2282 3088
rect 2226 3032 2228 3052
rect 2228 3032 2280 3052
rect 2280 3032 2282 3052
rect 3238 5072 3294 5128
rect 2930 4922 2986 4924
rect 3010 4922 3066 4924
rect 3090 4922 3146 4924
rect 3170 4922 3226 4924
rect 2930 4870 2976 4922
rect 2976 4870 2986 4922
rect 3010 4870 3040 4922
rect 3040 4870 3052 4922
rect 3052 4870 3066 4922
rect 3090 4870 3104 4922
rect 3104 4870 3116 4922
rect 3116 4870 3146 4922
rect 3170 4870 3180 4922
rect 3180 4870 3226 4922
rect 2930 4868 2986 4870
rect 3010 4868 3066 4870
rect 3090 4868 3146 4870
rect 3170 4868 3226 4870
rect 3054 4664 3110 4720
rect 2870 4140 2926 4176
rect 2870 4120 2872 4140
rect 2872 4120 2924 4140
rect 2924 4120 2926 4140
rect 2930 3834 2986 3836
rect 3010 3834 3066 3836
rect 3090 3834 3146 3836
rect 3170 3834 3226 3836
rect 2930 3782 2976 3834
rect 2976 3782 2986 3834
rect 3010 3782 3040 3834
rect 3040 3782 3052 3834
rect 3052 3782 3066 3834
rect 3090 3782 3104 3834
rect 3104 3782 3116 3834
rect 3116 3782 3146 3834
rect 3170 3782 3180 3834
rect 3180 3782 3226 3834
rect 2930 3780 2986 3782
rect 3010 3780 3066 3782
rect 3090 3780 3146 3782
rect 3170 3780 3226 3782
rect 2778 3576 2834 3632
rect 2962 3476 2964 3496
rect 2964 3476 3016 3496
rect 3016 3476 3018 3496
rect 2962 3440 3018 3476
rect 3146 3304 3202 3360
rect 4250 11600 4306 11656
rect 4710 15408 4766 15464
rect 4904 15258 4960 15260
rect 4984 15258 5040 15260
rect 5064 15258 5120 15260
rect 5144 15258 5200 15260
rect 4904 15206 4950 15258
rect 4950 15206 4960 15258
rect 4984 15206 5014 15258
rect 5014 15206 5026 15258
rect 5026 15206 5040 15258
rect 5064 15206 5078 15258
rect 5078 15206 5090 15258
rect 5090 15206 5120 15258
rect 5144 15206 5154 15258
rect 5154 15206 5200 15258
rect 4904 15204 4960 15206
rect 4984 15204 5040 15206
rect 5064 15204 5120 15206
rect 5144 15204 5200 15206
rect 4904 14170 4960 14172
rect 4984 14170 5040 14172
rect 5064 14170 5120 14172
rect 5144 14170 5200 14172
rect 4904 14118 4950 14170
rect 4950 14118 4960 14170
rect 4984 14118 5014 14170
rect 5014 14118 5026 14170
rect 5026 14118 5040 14170
rect 5064 14118 5078 14170
rect 5078 14118 5090 14170
rect 5090 14118 5120 14170
rect 5144 14118 5154 14170
rect 5154 14118 5200 14170
rect 4904 14116 4960 14118
rect 4984 14116 5040 14118
rect 5064 14116 5120 14118
rect 5144 14116 5200 14118
rect 5722 15564 5778 15600
rect 5722 15544 5724 15564
rect 5724 15544 5776 15564
rect 5776 15544 5778 15564
rect 5814 15408 5870 15464
rect 5446 14048 5502 14104
rect 5998 14320 6054 14376
rect 5722 13912 5778 13968
rect 4904 13082 4960 13084
rect 4984 13082 5040 13084
rect 5064 13082 5120 13084
rect 5144 13082 5200 13084
rect 4904 13030 4950 13082
rect 4950 13030 4960 13082
rect 4984 13030 5014 13082
rect 5014 13030 5026 13082
rect 5026 13030 5040 13082
rect 5064 13030 5078 13082
rect 5078 13030 5090 13082
rect 5090 13030 5120 13082
rect 5144 13030 5154 13082
rect 5154 13030 5200 13082
rect 4904 13028 4960 13030
rect 4984 13028 5040 13030
rect 5064 13028 5120 13030
rect 5144 13028 5200 13030
rect 4710 12824 4766 12880
rect 5538 12688 5594 12744
rect 4986 12552 5042 12608
rect 4904 11994 4960 11996
rect 4984 11994 5040 11996
rect 5064 11994 5120 11996
rect 5144 11994 5200 11996
rect 4904 11942 4950 11994
rect 4950 11942 4960 11994
rect 4984 11942 5014 11994
rect 5014 11942 5026 11994
rect 5026 11942 5040 11994
rect 5064 11942 5078 11994
rect 5078 11942 5090 11994
rect 5090 11942 5120 11994
rect 5144 11942 5154 11994
rect 5154 11942 5200 11994
rect 4904 11940 4960 11942
rect 4984 11940 5040 11942
rect 5064 11940 5120 11942
rect 5144 11940 5200 11942
rect 4904 10906 4960 10908
rect 4984 10906 5040 10908
rect 5064 10906 5120 10908
rect 5144 10906 5200 10908
rect 4904 10854 4950 10906
rect 4950 10854 4960 10906
rect 4984 10854 5014 10906
rect 5014 10854 5026 10906
rect 5026 10854 5040 10906
rect 5064 10854 5078 10906
rect 5078 10854 5090 10906
rect 5090 10854 5120 10906
rect 5144 10854 5154 10906
rect 5154 10854 5200 10906
rect 4904 10852 4960 10854
rect 4984 10852 5040 10854
rect 5064 10852 5120 10854
rect 5144 10852 5200 10854
rect 4066 9968 4122 10024
rect 3514 8916 3516 8936
rect 3516 8916 3568 8936
rect 3568 8916 3570 8936
rect 3514 8880 3570 8916
rect 3514 8336 3570 8392
rect 3422 7928 3478 7984
rect 2930 2746 2986 2748
rect 3010 2746 3066 2748
rect 3090 2746 3146 2748
rect 3170 2746 3226 2748
rect 2930 2694 2976 2746
rect 2976 2694 2986 2746
rect 3010 2694 3040 2746
rect 3040 2694 3052 2746
rect 3052 2694 3066 2746
rect 3090 2694 3104 2746
rect 3104 2694 3116 2746
rect 3116 2694 3146 2746
rect 3170 2694 3180 2746
rect 3180 2694 3226 2746
rect 2930 2692 2986 2694
rect 3010 2692 3066 2694
rect 3090 2692 3146 2694
rect 3170 2692 3226 2694
rect 3606 4256 3662 4312
rect 3974 8200 4030 8256
rect 3882 6024 3938 6080
rect 4250 7384 4306 7440
rect 4158 6976 4214 7032
rect 4066 6860 4122 6896
rect 4066 6840 4068 6860
rect 4068 6840 4120 6860
rect 4120 6840 4122 6860
rect 3974 5752 4030 5808
rect 3790 5208 3846 5264
rect 3974 5228 4030 5264
rect 3974 5208 3976 5228
rect 3976 5208 4028 5228
rect 4028 5208 4030 5228
rect 4066 4820 4122 4856
rect 4066 4800 4068 4820
rect 4068 4800 4120 4820
rect 4120 4800 4122 4820
rect 3974 4020 3976 4040
rect 3976 4020 4028 4040
rect 4028 4020 4030 4040
rect 3974 3984 4030 4020
rect 4904 9818 4960 9820
rect 4984 9818 5040 9820
rect 5064 9818 5120 9820
rect 5144 9818 5200 9820
rect 4904 9766 4950 9818
rect 4950 9766 4960 9818
rect 4984 9766 5014 9818
rect 5014 9766 5026 9818
rect 5026 9766 5040 9818
rect 5064 9766 5078 9818
rect 5078 9766 5090 9818
rect 5090 9766 5120 9818
rect 5144 9766 5154 9818
rect 5154 9766 5200 9818
rect 4904 9764 4960 9766
rect 4984 9764 5040 9766
rect 5064 9764 5120 9766
rect 5144 9764 5200 9766
rect 4710 8472 4766 8528
rect 4710 7928 4766 7984
rect 4710 6704 4766 6760
rect 4904 8730 4960 8732
rect 4984 8730 5040 8732
rect 5064 8730 5120 8732
rect 5144 8730 5200 8732
rect 4904 8678 4950 8730
rect 4950 8678 4960 8730
rect 4984 8678 5014 8730
rect 5014 8678 5026 8730
rect 5026 8678 5040 8730
rect 5064 8678 5078 8730
rect 5078 8678 5090 8730
rect 5090 8678 5120 8730
rect 5144 8678 5154 8730
rect 5154 8678 5200 8730
rect 4904 8676 4960 8678
rect 4984 8676 5040 8678
rect 5064 8676 5120 8678
rect 5144 8676 5200 8678
rect 5078 8472 5134 8528
rect 4904 7642 4960 7644
rect 4984 7642 5040 7644
rect 5064 7642 5120 7644
rect 5144 7642 5200 7644
rect 4904 7590 4950 7642
rect 4950 7590 4960 7642
rect 4984 7590 5014 7642
rect 5014 7590 5026 7642
rect 5026 7590 5040 7642
rect 5064 7590 5078 7642
rect 5078 7590 5090 7642
rect 5090 7590 5120 7642
rect 5144 7590 5154 7642
rect 5154 7590 5200 7642
rect 4904 7588 4960 7590
rect 4984 7588 5040 7590
rect 5064 7588 5120 7590
rect 5144 7588 5200 7590
rect 5170 6996 5226 7032
rect 5170 6976 5172 6996
rect 5172 6976 5224 6996
rect 5224 6976 5226 6996
rect 4904 6554 4960 6556
rect 4984 6554 5040 6556
rect 5064 6554 5120 6556
rect 5144 6554 5200 6556
rect 4904 6502 4950 6554
rect 4950 6502 4960 6554
rect 4984 6502 5014 6554
rect 5014 6502 5026 6554
rect 5026 6502 5040 6554
rect 5064 6502 5078 6554
rect 5078 6502 5090 6554
rect 5090 6502 5120 6554
rect 5144 6502 5154 6554
rect 5154 6502 5200 6554
rect 4904 6500 4960 6502
rect 4984 6500 5040 6502
rect 5064 6500 5120 6502
rect 5144 6500 5200 6502
rect 4986 5752 5042 5808
rect 5078 5616 5134 5672
rect 4904 5466 4960 5468
rect 4984 5466 5040 5468
rect 5064 5466 5120 5468
rect 5144 5466 5200 5468
rect 4904 5414 4950 5466
rect 4950 5414 4960 5466
rect 4984 5414 5014 5466
rect 5014 5414 5026 5466
rect 5026 5414 5040 5466
rect 5064 5414 5078 5466
rect 5078 5414 5090 5466
rect 5090 5414 5120 5466
rect 5144 5414 5154 5466
rect 5154 5414 5200 5466
rect 4904 5412 4960 5414
rect 4984 5412 5040 5414
rect 5064 5412 5120 5414
rect 5144 5412 5200 5414
rect 4710 4972 4712 4992
rect 4712 4972 4764 4992
rect 4764 4972 4766 4992
rect 4710 4936 4766 4972
rect 4904 4378 4960 4380
rect 4984 4378 5040 4380
rect 5064 4378 5120 4380
rect 5144 4378 5200 4380
rect 4904 4326 4950 4378
rect 4950 4326 4960 4378
rect 4984 4326 5014 4378
rect 5014 4326 5026 4378
rect 5026 4326 5040 4378
rect 5064 4326 5078 4378
rect 5078 4326 5090 4378
rect 5090 4326 5120 4378
rect 5144 4326 5154 4378
rect 5154 4326 5200 4378
rect 4904 4324 4960 4326
rect 4984 4324 5040 4326
rect 5064 4324 5120 4326
rect 5144 4324 5200 4326
rect 5630 10648 5686 10704
rect 6878 16890 6934 16892
rect 6958 16890 7014 16892
rect 7038 16890 7094 16892
rect 7118 16890 7174 16892
rect 6878 16838 6924 16890
rect 6924 16838 6934 16890
rect 6958 16838 6988 16890
rect 6988 16838 7000 16890
rect 7000 16838 7014 16890
rect 7038 16838 7052 16890
rect 7052 16838 7064 16890
rect 7064 16838 7094 16890
rect 7118 16838 7128 16890
rect 7128 16838 7174 16890
rect 6878 16836 6934 16838
rect 6958 16836 7014 16838
rect 7038 16836 7094 16838
rect 7118 16836 7174 16838
rect 10826 16890 10882 16892
rect 10906 16890 10962 16892
rect 10986 16890 11042 16892
rect 11066 16890 11122 16892
rect 10826 16838 10872 16890
rect 10872 16838 10882 16890
rect 10906 16838 10936 16890
rect 10936 16838 10948 16890
rect 10948 16838 10962 16890
rect 10986 16838 11000 16890
rect 11000 16838 11012 16890
rect 11012 16838 11042 16890
rect 11066 16838 11076 16890
rect 11076 16838 11122 16890
rect 10826 16836 10882 16838
rect 10906 16836 10962 16838
rect 10986 16836 11042 16838
rect 11066 16836 11122 16838
rect 6366 14884 6422 14920
rect 6366 14864 6368 14884
rect 6368 14864 6420 14884
rect 6420 14864 6422 14884
rect 5722 8064 5778 8120
rect 8852 16346 8908 16348
rect 8932 16346 8988 16348
rect 9012 16346 9068 16348
rect 9092 16346 9148 16348
rect 8852 16294 8898 16346
rect 8898 16294 8908 16346
rect 8932 16294 8962 16346
rect 8962 16294 8974 16346
rect 8974 16294 8988 16346
rect 9012 16294 9026 16346
rect 9026 16294 9038 16346
rect 9038 16294 9068 16346
rect 9092 16294 9102 16346
rect 9102 16294 9148 16346
rect 8852 16292 8908 16294
rect 8932 16292 8988 16294
rect 9012 16292 9068 16294
rect 9092 16292 9148 16294
rect 6878 15802 6934 15804
rect 6958 15802 7014 15804
rect 7038 15802 7094 15804
rect 7118 15802 7174 15804
rect 6878 15750 6924 15802
rect 6924 15750 6934 15802
rect 6958 15750 6988 15802
rect 6988 15750 7000 15802
rect 7000 15750 7014 15802
rect 7038 15750 7052 15802
rect 7052 15750 7064 15802
rect 7064 15750 7094 15802
rect 7118 15750 7128 15802
rect 7128 15750 7174 15802
rect 6878 15748 6934 15750
rect 6958 15748 7014 15750
rect 7038 15748 7094 15750
rect 7118 15748 7174 15750
rect 7102 14864 7158 14920
rect 6878 14714 6934 14716
rect 6958 14714 7014 14716
rect 7038 14714 7094 14716
rect 7118 14714 7174 14716
rect 6878 14662 6924 14714
rect 6924 14662 6934 14714
rect 6958 14662 6988 14714
rect 6988 14662 7000 14714
rect 7000 14662 7014 14714
rect 7038 14662 7052 14714
rect 7052 14662 7064 14714
rect 7064 14662 7094 14714
rect 7118 14662 7128 14714
rect 7128 14662 7174 14714
rect 6878 14660 6934 14662
rect 6958 14660 7014 14662
rect 7038 14660 7094 14662
rect 7118 14660 7174 14662
rect 6878 13626 6934 13628
rect 6958 13626 7014 13628
rect 7038 13626 7094 13628
rect 7118 13626 7174 13628
rect 6878 13574 6924 13626
rect 6924 13574 6934 13626
rect 6958 13574 6988 13626
rect 6988 13574 7000 13626
rect 7000 13574 7014 13626
rect 7038 13574 7052 13626
rect 7052 13574 7064 13626
rect 7064 13574 7094 13626
rect 7118 13574 7128 13626
rect 7128 13574 7174 13626
rect 6878 13572 6934 13574
rect 6958 13572 7014 13574
rect 7038 13572 7094 13574
rect 7118 13572 7174 13574
rect 6734 13368 6790 13424
rect 6878 12538 6934 12540
rect 6958 12538 7014 12540
rect 7038 12538 7094 12540
rect 7118 12538 7174 12540
rect 6878 12486 6924 12538
rect 6924 12486 6934 12538
rect 6958 12486 6988 12538
rect 6988 12486 7000 12538
rect 7000 12486 7014 12538
rect 7038 12486 7052 12538
rect 7052 12486 7064 12538
rect 7064 12486 7094 12538
rect 7118 12486 7128 12538
rect 7128 12486 7174 12538
rect 6878 12484 6934 12486
rect 6958 12484 7014 12486
rect 7038 12484 7094 12486
rect 7118 12484 7174 12486
rect 6734 12280 6790 12336
rect 6642 11464 6698 11520
rect 6090 8916 6092 8936
rect 6092 8916 6144 8936
rect 6144 8916 6146 8936
rect 6090 8880 6146 8916
rect 6182 8064 6238 8120
rect 6366 8064 6422 8120
rect 5538 7656 5594 7712
rect 5906 7520 5962 7576
rect 6366 7928 6422 7984
rect 6550 9016 6606 9072
rect 5630 7112 5686 7168
rect 5630 6840 5686 6896
rect 5446 5616 5502 5672
rect 5354 5364 5410 5400
rect 5354 5344 5356 5364
rect 5356 5344 5408 5364
rect 5408 5344 5410 5364
rect 5630 5344 5686 5400
rect 5814 6568 5870 6624
rect 5814 5480 5870 5536
rect 6826 12144 6882 12200
rect 6878 11450 6934 11452
rect 6958 11450 7014 11452
rect 7038 11450 7094 11452
rect 7118 11450 7174 11452
rect 6878 11398 6924 11450
rect 6924 11398 6934 11450
rect 6958 11398 6988 11450
rect 6988 11398 7000 11450
rect 7000 11398 7014 11450
rect 7038 11398 7052 11450
rect 7052 11398 7064 11450
rect 7064 11398 7094 11450
rect 7118 11398 7128 11450
rect 7128 11398 7174 11450
rect 6878 11396 6934 11398
rect 6958 11396 7014 11398
rect 7038 11396 7094 11398
rect 7118 11396 7174 11398
rect 6878 10362 6934 10364
rect 6958 10362 7014 10364
rect 7038 10362 7094 10364
rect 7118 10362 7174 10364
rect 6878 10310 6924 10362
rect 6924 10310 6934 10362
rect 6958 10310 6988 10362
rect 6988 10310 7000 10362
rect 7000 10310 7014 10362
rect 7038 10310 7052 10362
rect 7052 10310 7064 10362
rect 7064 10310 7094 10362
rect 7118 10310 7128 10362
rect 7128 10310 7174 10362
rect 6878 10308 6934 10310
rect 6958 10308 7014 10310
rect 7038 10308 7094 10310
rect 7118 10308 7174 10310
rect 7654 15000 7710 15056
rect 7562 14048 7618 14104
rect 7470 11600 7526 11656
rect 6878 9274 6934 9276
rect 6958 9274 7014 9276
rect 7038 9274 7094 9276
rect 7118 9274 7174 9276
rect 6878 9222 6924 9274
rect 6924 9222 6934 9274
rect 6958 9222 6988 9274
rect 6988 9222 7000 9274
rect 7000 9222 7014 9274
rect 7038 9222 7052 9274
rect 7052 9222 7064 9274
rect 7064 9222 7094 9274
rect 7118 9222 7128 9274
rect 7128 9222 7174 9274
rect 6878 9220 6934 9222
rect 6958 9220 7014 9222
rect 7038 9220 7094 9222
rect 7118 9220 7174 9222
rect 7102 8880 7158 8936
rect 6826 8472 6882 8528
rect 6878 8186 6934 8188
rect 6958 8186 7014 8188
rect 7038 8186 7094 8188
rect 7118 8186 7174 8188
rect 6878 8134 6924 8186
rect 6924 8134 6934 8186
rect 6958 8134 6988 8186
rect 6988 8134 7000 8186
rect 7000 8134 7014 8186
rect 7038 8134 7052 8186
rect 7052 8134 7064 8186
rect 7064 8134 7094 8186
rect 7118 8134 7128 8186
rect 7128 8134 7174 8186
rect 6878 8132 6934 8134
rect 6958 8132 7014 8134
rect 7038 8132 7094 8134
rect 7118 8132 7174 8134
rect 7102 7964 7104 7984
rect 7104 7964 7156 7984
rect 7156 7964 7158 7984
rect 7102 7928 7158 7964
rect 7102 7520 7158 7576
rect 6826 7384 6882 7440
rect 6366 7112 6422 7168
rect 6366 6840 6422 6896
rect 6090 6568 6146 6624
rect 6182 6432 6238 6488
rect 6550 6432 6606 6488
rect 6550 6024 6606 6080
rect 6182 4820 6238 4856
rect 6182 4800 6184 4820
rect 6184 4800 6236 4820
rect 6236 4800 6238 4820
rect 6878 7098 6934 7100
rect 6958 7098 7014 7100
rect 7038 7098 7094 7100
rect 7118 7098 7174 7100
rect 6878 7046 6924 7098
rect 6924 7046 6934 7098
rect 6958 7046 6988 7098
rect 6988 7046 7000 7098
rect 7000 7046 7014 7098
rect 7038 7046 7052 7098
rect 7052 7046 7064 7098
rect 7064 7046 7094 7098
rect 7118 7046 7128 7098
rect 7128 7046 7174 7098
rect 6878 7044 6934 7046
rect 6958 7044 7014 7046
rect 7038 7044 7094 7046
rect 7118 7044 7174 7046
rect 6918 6432 6974 6488
rect 7286 6840 7342 6896
rect 6878 6010 6934 6012
rect 6958 6010 7014 6012
rect 7038 6010 7094 6012
rect 7118 6010 7174 6012
rect 6878 5958 6924 6010
rect 6924 5958 6934 6010
rect 6958 5958 6988 6010
rect 6988 5958 7000 6010
rect 7000 5958 7014 6010
rect 7038 5958 7052 6010
rect 7052 5958 7064 6010
rect 7064 5958 7094 6010
rect 7118 5958 7128 6010
rect 7128 5958 7174 6010
rect 6878 5956 6934 5958
rect 6958 5956 7014 5958
rect 7038 5956 7094 5958
rect 7118 5956 7174 5958
rect 7654 10240 7710 10296
rect 8852 15258 8908 15260
rect 8932 15258 8988 15260
rect 9012 15258 9068 15260
rect 9092 15258 9148 15260
rect 8852 15206 8898 15258
rect 8898 15206 8908 15258
rect 8932 15206 8962 15258
rect 8962 15206 8974 15258
rect 8974 15206 8988 15258
rect 9012 15206 9026 15258
rect 9026 15206 9038 15258
rect 9038 15206 9068 15258
rect 9092 15206 9102 15258
rect 9102 15206 9148 15258
rect 8852 15204 8908 15206
rect 8932 15204 8988 15206
rect 9012 15204 9068 15206
rect 9092 15204 9148 15206
rect 8022 13368 8078 13424
rect 8114 12824 8170 12880
rect 8022 12552 8078 12608
rect 7930 11736 7986 11792
rect 8852 14170 8908 14172
rect 8932 14170 8988 14172
rect 9012 14170 9068 14172
rect 9092 14170 9148 14172
rect 8852 14118 8898 14170
rect 8898 14118 8908 14170
rect 8932 14118 8962 14170
rect 8962 14118 8974 14170
rect 8974 14118 8988 14170
rect 9012 14118 9026 14170
rect 9026 14118 9038 14170
rect 9038 14118 9068 14170
rect 9092 14118 9102 14170
rect 9102 14118 9148 14170
rect 8852 14116 8908 14118
rect 8932 14116 8988 14118
rect 9012 14116 9068 14118
rect 9092 14116 9148 14118
rect 8666 13232 8722 13288
rect 8852 13082 8908 13084
rect 8932 13082 8988 13084
rect 9012 13082 9068 13084
rect 9092 13082 9148 13084
rect 8852 13030 8898 13082
rect 8898 13030 8908 13082
rect 8932 13030 8962 13082
rect 8962 13030 8974 13082
rect 8974 13030 8988 13082
rect 9012 13030 9026 13082
rect 9026 13030 9038 13082
rect 9038 13030 9068 13082
rect 9092 13030 9102 13082
rect 9102 13030 9148 13082
rect 8852 13028 8908 13030
rect 8932 13028 8988 13030
rect 9012 13028 9068 13030
rect 9092 13028 9148 13030
rect 7838 11600 7894 11656
rect 7838 11192 7894 11248
rect 7654 9288 7710 9344
rect 7654 9152 7710 9208
rect 8206 11736 8262 11792
rect 7562 8356 7618 8392
rect 7562 8336 7564 8356
rect 7564 8336 7616 8356
rect 7616 8336 7618 8356
rect 8022 9016 8078 9072
rect 7470 7792 7526 7848
rect 7562 6860 7618 6896
rect 7562 6840 7564 6860
rect 7564 6840 7616 6860
rect 7616 6840 7618 6860
rect 7562 5616 7618 5672
rect 6878 4922 6934 4924
rect 6958 4922 7014 4924
rect 7038 4922 7094 4924
rect 7118 4922 7174 4924
rect 6878 4870 6924 4922
rect 6924 4870 6934 4922
rect 6958 4870 6988 4922
rect 6988 4870 7000 4922
rect 7000 4870 7014 4922
rect 7038 4870 7052 4922
rect 7052 4870 7064 4922
rect 7064 4870 7094 4922
rect 7118 4870 7128 4922
rect 7128 4870 7174 4922
rect 6878 4868 6934 4870
rect 6958 4868 7014 4870
rect 7038 4868 7094 4870
rect 7118 4868 7174 4870
rect 6642 4564 6644 4584
rect 6644 4564 6696 4584
rect 6696 4564 6698 4584
rect 5722 4120 5778 4176
rect 6642 4528 6698 4564
rect 5630 3848 5686 3904
rect 4904 3290 4960 3292
rect 4984 3290 5040 3292
rect 5064 3290 5120 3292
rect 5144 3290 5200 3292
rect 4904 3238 4950 3290
rect 4950 3238 4960 3290
rect 4984 3238 5014 3290
rect 5014 3238 5026 3290
rect 5026 3238 5040 3290
rect 5064 3238 5078 3290
rect 5078 3238 5090 3290
rect 5090 3238 5120 3290
rect 5144 3238 5154 3290
rect 5154 3238 5200 3290
rect 4904 3236 4960 3238
rect 4984 3236 5040 3238
rect 5064 3236 5120 3238
rect 5144 3236 5200 3238
rect 7286 4120 7342 4176
rect 8206 9444 8262 9480
rect 8206 9424 8208 9444
rect 8208 9424 8260 9444
rect 8260 9424 8262 9444
rect 8206 9288 8262 9344
rect 8206 8744 8262 8800
rect 7838 7520 7894 7576
rect 7838 7112 7894 7168
rect 7838 5652 7840 5672
rect 7840 5652 7892 5672
rect 7892 5652 7894 5672
rect 7654 5344 7710 5400
rect 7838 5616 7894 5652
rect 6878 3834 6934 3836
rect 6958 3834 7014 3836
rect 7038 3834 7094 3836
rect 7118 3834 7174 3836
rect 6878 3782 6924 3834
rect 6924 3782 6934 3834
rect 6958 3782 6988 3834
rect 6988 3782 7000 3834
rect 7000 3782 7014 3834
rect 7038 3782 7052 3834
rect 7052 3782 7064 3834
rect 7064 3782 7094 3834
rect 7118 3782 7128 3834
rect 7128 3782 7174 3834
rect 6878 3780 6934 3782
rect 6958 3780 7014 3782
rect 7038 3780 7094 3782
rect 7118 3780 7174 3782
rect 8574 12008 8630 12064
rect 9034 12688 9090 12744
rect 8850 12416 8906 12472
rect 10826 15802 10882 15804
rect 10906 15802 10962 15804
rect 10986 15802 11042 15804
rect 11066 15802 11122 15804
rect 10826 15750 10872 15802
rect 10872 15750 10882 15802
rect 10906 15750 10936 15802
rect 10936 15750 10948 15802
rect 10948 15750 10962 15802
rect 10986 15750 11000 15802
rect 11000 15750 11012 15802
rect 11012 15750 11042 15802
rect 11066 15750 11076 15802
rect 11076 15750 11122 15802
rect 10826 15748 10882 15750
rect 10906 15748 10962 15750
rect 10986 15748 11042 15750
rect 11066 15748 11122 15750
rect 9126 12280 9182 12336
rect 10826 14714 10882 14716
rect 10906 14714 10962 14716
rect 10986 14714 11042 14716
rect 11066 14714 11122 14716
rect 10826 14662 10872 14714
rect 10872 14662 10882 14714
rect 10906 14662 10936 14714
rect 10936 14662 10948 14714
rect 10948 14662 10962 14714
rect 10986 14662 11000 14714
rect 11000 14662 11012 14714
rect 11012 14662 11042 14714
rect 11066 14662 11076 14714
rect 11076 14662 11122 14714
rect 10826 14660 10882 14662
rect 10906 14660 10962 14662
rect 10986 14660 11042 14662
rect 11066 14660 11122 14662
rect 10598 14320 10654 14376
rect 10322 13912 10378 13968
rect 9494 12416 9550 12472
rect 8852 11994 8908 11996
rect 8932 11994 8988 11996
rect 9012 11994 9068 11996
rect 9092 11994 9148 11996
rect 8852 11942 8898 11994
rect 8898 11942 8908 11994
rect 8932 11942 8962 11994
rect 8962 11942 8974 11994
rect 8974 11942 8988 11994
rect 9012 11942 9026 11994
rect 9026 11942 9038 11994
rect 9038 11942 9068 11994
rect 9092 11942 9102 11994
rect 9102 11942 9148 11994
rect 8852 11940 8908 11942
rect 8932 11940 8988 11942
rect 9012 11940 9068 11942
rect 9092 11940 9148 11942
rect 8850 11192 8906 11248
rect 9678 12280 9734 12336
rect 9586 12008 9642 12064
rect 9402 11756 9458 11792
rect 9402 11736 9404 11756
rect 9404 11736 9456 11756
rect 9456 11736 9458 11756
rect 9126 11464 9182 11520
rect 9034 11056 9090 11112
rect 9218 11056 9274 11112
rect 8852 10906 8908 10908
rect 8932 10906 8988 10908
rect 9012 10906 9068 10908
rect 9092 10906 9148 10908
rect 8852 10854 8898 10906
rect 8898 10854 8908 10906
rect 8932 10854 8962 10906
rect 8962 10854 8974 10906
rect 8974 10854 8988 10906
rect 9012 10854 9026 10906
rect 9026 10854 9038 10906
rect 9038 10854 9068 10906
rect 9092 10854 9102 10906
rect 9102 10854 9148 10906
rect 8852 10852 8908 10854
rect 8932 10852 8988 10854
rect 9012 10852 9068 10854
rect 9092 10852 9148 10854
rect 8758 10648 8814 10704
rect 8942 10648 8998 10704
rect 8942 10240 8998 10296
rect 9678 11464 9734 11520
rect 8852 9818 8908 9820
rect 8932 9818 8988 9820
rect 9012 9818 9068 9820
rect 9092 9818 9148 9820
rect 8852 9766 8898 9818
rect 8898 9766 8908 9818
rect 8932 9766 8962 9818
rect 8962 9766 8974 9818
rect 8974 9766 8988 9818
rect 9012 9766 9026 9818
rect 9026 9766 9038 9818
rect 9038 9766 9068 9818
rect 9092 9766 9102 9818
rect 9102 9766 9148 9818
rect 8852 9764 8908 9766
rect 8932 9764 8988 9766
rect 9012 9764 9068 9766
rect 9092 9764 9148 9766
rect 8574 9288 8630 9344
rect 8666 9016 8722 9072
rect 8574 8608 8630 8664
rect 8390 7656 8446 7712
rect 8482 6296 8538 6352
rect 9402 9324 9404 9344
rect 9404 9324 9456 9344
rect 9456 9324 9458 9344
rect 9402 9288 9458 9324
rect 8852 8730 8908 8732
rect 8932 8730 8988 8732
rect 9012 8730 9068 8732
rect 9092 8730 9148 8732
rect 8852 8678 8898 8730
rect 8898 8678 8908 8730
rect 8932 8678 8962 8730
rect 8962 8678 8974 8730
rect 8974 8678 8988 8730
rect 9012 8678 9026 8730
rect 9026 8678 9038 8730
rect 9038 8678 9068 8730
rect 9092 8678 9102 8730
rect 9102 8678 9148 8730
rect 8852 8676 8908 8678
rect 8932 8676 8988 8678
rect 9012 8676 9068 8678
rect 9092 8676 9148 8678
rect 9034 8336 9090 8392
rect 8942 8064 8998 8120
rect 8852 7642 8908 7644
rect 8932 7642 8988 7644
rect 9012 7642 9068 7644
rect 9092 7642 9148 7644
rect 8852 7590 8898 7642
rect 8898 7590 8908 7642
rect 8932 7590 8962 7642
rect 8962 7590 8974 7642
rect 8974 7590 8988 7642
rect 9012 7590 9026 7642
rect 9026 7590 9038 7642
rect 9038 7590 9068 7642
rect 9092 7590 9102 7642
rect 9102 7590 9148 7642
rect 8852 7588 8908 7590
rect 8932 7588 8988 7590
rect 9012 7588 9068 7590
rect 9092 7588 9148 7590
rect 9034 7384 9090 7440
rect 9678 10804 9734 10840
rect 10138 12824 10194 12880
rect 10138 11600 10194 11656
rect 10138 11192 10194 11248
rect 9678 10784 9680 10804
rect 9680 10784 9732 10804
rect 9732 10784 9734 10804
rect 9862 10376 9918 10432
rect 9586 9832 9642 9888
rect 9678 9152 9734 9208
rect 10046 9696 10102 9752
rect 9954 9424 10010 9480
rect 10506 11464 10562 11520
rect 10826 13626 10882 13628
rect 10906 13626 10962 13628
rect 10986 13626 11042 13628
rect 11066 13626 11122 13628
rect 10826 13574 10872 13626
rect 10872 13574 10882 13626
rect 10906 13574 10936 13626
rect 10936 13574 10948 13626
rect 10948 13574 10962 13626
rect 10986 13574 11000 13626
rect 11000 13574 11012 13626
rect 11012 13574 11042 13626
rect 11066 13574 11076 13626
rect 11076 13574 11122 13626
rect 10826 13572 10882 13574
rect 10906 13572 10962 13574
rect 10986 13572 11042 13574
rect 11066 13572 11122 13574
rect 10826 12538 10882 12540
rect 10906 12538 10962 12540
rect 10986 12538 11042 12540
rect 11066 12538 11122 12540
rect 10826 12486 10872 12538
rect 10872 12486 10882 12538
rect 10906 12486 10936 12538
rect 10936 12486 10948 12538
rect 10948 12486 10962 12538
rect 10986 12486 11000 12538
rect 11000 12486 11012 12538
rect 11012 12486 11042 12538
rect 11066 12486 11076 12538
rect 11076 12486 11122 12538
rect 10826 12484 10882 12486
rect 10906 12484 10962 12486
rect 10986 12484 11042 12486
rect 11066 12484 11122 12486
rect 10782 12280 10838 12336
rect 10690 11736 10746 11792
rect 10826 11450 10882 11452
rect 10906 11450 10962 11452
rect 10986 11450 11042 11452
rect 11066 11450 11122 11452
rect 10826 11398 10872 11450
rect 10872 11398 10882 11450
rect 10906 11398 10936 11450
rect 10936 11398 10948 11450
rect 10948 11398 10962 11450
rect 10986 11398 11000 11450
rect 11000 11398 11012 11450
rect 11012 11398 11042 11450
rect 11066 11398 11076 11450
rect 11076 11398 11122 11450
rect 10826 11396 10882 11398
rect 10906 11396 10962 11398
rect 10986 11396 11042 11398
rect 11066 11396 11122 11398
rect 11150 11192 11206 11248
rect 10782 11076 10838 11112
rect 10782 11056 10784 11076
rect 10784 11056 10836 11076
rect 10836 11056 10838 11076
rect 14774 16890 14830 16892
rect 14854 16890 14910 16892
rect 14934 16890 14990 16892
rect 15014 16890 15070 16892
rect 14774 16838 14820 16890
rect 14820 16838 14830 16890
rect 14854 16838 14884 16890
rect 14884 16838 14896 16890
rect 14896 16838 14910 16890
rect 14934 16838 14948 16890
rect 14948 16838 14960 16890
rect 14960 16838 14990 16890
rect 15014 16838 15024 16890
rect 15024 16838 15070 16890
rect 14774 16836 14830 16838
rect 14854 16836 14910 16838
rect 14934 16836 14990 16838
rect 15014 16836 15070 16838
rect 12800 16346 12856 16348
rect 12880 16346 12936 16348
rect 12960 16346 13016 16348
rect 13040 16346 13096 16348
rect 12800 16294 12846 16346
rect 12846 16294 12856 16346
rect 12880 16294 12910 16346
rect 12910 16294 12922 16346
rect 12922 16294 12936 16346
rect 12960 16294 12974 16346
rect 12974 16294 12986 16346
rect 12986 16294 13016 16346
rect 13040 16294 13050 16346
rect 13050 16294 13096 16346
rect 12800 16292 12856 16294
rect 12880 16292 12936 16294
rect 12960 16292 13016 16294
rect 13040 16292 13096 16294
rect 14774 15802 14830 15804
rect 14854 15802 14910 15804
rect 14934 15802 14990 15804
rect 15014 15802 15070 15804
rect 14774 15750 14820 15802
rect 14820 15750 14830 15802
rect 14854 15750 14884 15802
rect 14884 15750 14896 15802
rect 14896 15750 14910 15802
rect 14934 15750 14948 15802
rect 14948 15750 14960 15802
rect 14960 15750 14990 15802
rect 15014 15750 15024 15802
rect 15024 15750 15070 15802
rect 14774 15748 14830 15750
rect 14854 15748 14910 15750
rect 14934 15748 14990 15750
rect 15014 15748 15070 15750
rect 12800 15258 12856 15260
rect 12880 15258 12936 15260
rect 12960 15258 13016 15260
rect 13040 15258 13096 15260
rect 12800 15206 12846 15258
rect 12846 15206 12856 15258
rect 12880 15206 12910 15258
rect 12910 15206 12922 15258
rect 12922 15206 12936 15258
rect 12960 15206 12974 15258
rect 12974 15206 12986 15258
rect 12986 15206 13016 15258
rect 13040 15206 13050 15258
rect 13050 15206 13096 15258
rect 12800 15204 12856 15206
rect 12880 15204 12936 15206
rect 12960 15204 13016 15206
rect 13040 15204 13096 15206
rect 14774 14714 14830 14716
rect 14854 14714 14910 14716
rect 14934 14714 14990 14716
rect 15014 14714 15070 14716
rect 14774 14662 14820 14714
rect 14820 14662 14830 14714
rect 14854 14662 14884 14714
rect 14884 14662 14896 14714
rect 14896 14662 14910 14714
rect 14934 14662 14948 14714
rect 14948 14662 14960 14714
rect 14960 14662 14990 14714
rect 15014 14662 15024 14714
rect 15024 14662 15070 14714
rect 14774 14660 14830 14662
rect 14854 14660 14910 14662
rect 14934 14660 14990 14662
rect 15014 14660 15070 14662
rect 12800 14170 12856 14172
rect 12880 14170 12936 14172
rect 12960 14170 13016 14172
rect 13040 14170 13096 14172
rect 12800 14118 12846 14170
rect 12846 14118 12856 14170
rect 12880 14118 12910 14170
rect 12910 14118 12922 14170
rect 12922 14118 12936 14170
rect 12960 14118 12974 14170
rect 12974 14118 12986 14170
rect 12986 14118 13016 14170
rect 13040 14118 13050 14170
rect 13050 14118 13096 14170
rect 12800 14116 12856 14118
rect 12880 14116 12936 14118
rect 12960 14116 13016 14118
rect 13040 14116 13096 14118
rect 10874 10784 10930 10840
rect 11150 10512 11206 10568
rect 10826 10362 10882 10364
rect 10906 10362 10962 10364
rect 10986 10362 11042 10364
rect 11066 10362 11122 10364
rect 10826 10310 10872 10362
rect 10872 10310 10882 10362
rect 10906 10310 10936 10362
rect 10936 10310 10948 10362
rect 10948 10310 10962 10362
rect 10986 10310 11000 10362
rect 11000 10310 11012 10362
rect 11012 10310 11042 10362
rect 11066 10310 11076 10362
rect 11076 10310 11122 10362
rect 10826 10308 10882 10310
rect 10906 10308 10962 10310
rect 10986 10308 11042 10310
rect 11066 10308 11122 10310
rect 10690 10240 10746 10296
rect 9862 9016 9918 9072
rect 10138 9288 10194 9344
rect 9402 7248 9458 7304
rect 9402 7148 9404 7168
rect 9404 7148 9456 7168
rect 9456 7148 9458 7168
rect 9402 7112 9458 7148
rect 8852 6554 8908 6556
rect 8932 6554 8988 6556
rect 9012 6554 9068 6556
rect 9092 6554 9148 6556
rect 8852 6502 8898 6554
rect 8898 6502 8908 6554
rect 8932 6502 8962 6554
rect 8962 6502 8974 6554
rect 8974 6502 8988 6554
rect 9012 6502 9026 6554
rect 9026 6502 9038 6554
rect 9038 6502 9068 6554
rect 9092 6502 9102 6554
rect 9102 6502 9148 6554
rect 8852 6500 8908 6502
rect 8932 6500 8988 6502
rect 9012 6500 9068 6502
rect 9092 6500 9148 6502
rect 8758 6296 8814 6352
rect 8758 6180 8814 6216
rect 8758 6160 8760 6180
rect 8760 6160 8812 6180
rect 8812 6160 8814 6180
rect 8852 5466 8908 5468
rect 8932 5466 8988 5468
rect 9012 5466 9068 5468
rect 9092 5466 9148 5468
rect 8852 5414 8898 5466
rect 8898 5414 8908 5466
rect 8932 5414 8962 5466
rect 8962 5414 8974 5466
rect 8974 5414 8988 5466
rect 9012 5414 9026 5466
rect 9026 5414 9038 5466
rect 9038 5414 9068 5466
rect 9092 5414 9102 5466
rect 9102 5414 9148 5466
rect 8852 5412 8908 5414
rect 8932 5412 8988 5414
rect 9012 5412 9068 5414
rect 9092 5412 9148 5414
rect 8482 5344 8538 5400
rect 10046 8336 10102 8392
rect 9678 7656 9734 7712
rect 9862 7520 9918 7576
rect 8852 4378 8908 4380
rect 8932 4378 8988 4380
rect 9012 4378 9068 4380
rect 9092 4378 9148 4380
rect 8852 4326 8898 4378
rect 8898 4326 8908 4378
rect 8932 4326 8962 4378
rect 8962 4326 8974 4378
rect 8974 4326 8988 4378
rect 9012 4326 9026 4378
rect 9026 4326 9038 4378
rect 9038 4326 9068 4378
rect 9092 4326 9102 4378
rect 9102 4326 9148 4378
rect 8852 4324 8908 4326
rect 8932 4324 8988 4326
rect 9012 4324 9068 4326
rect 9092 4324 9148 4326
rect 8852 3290 8908 3292
rect 8932 3290 8988 3292
rect 9012 3290 9068 3292
rect 9092 3290 9148 3292
rect 8852 3238 8898 3290
rect 8898 3238 8908 3290
rect 8932 3238 8962 3290
rect 8962 3238 8974 3290
rect 8974 3238 8988 3290
rect 9012 3238 9026 3290
rect 9026 3238 9038 3290
rect 9038 3238 9068 3290
rect 9092 3238 9102 3290
rect 9102 3238 9148 3290
rect 8852 3236 8908 3238
rect 8932 3236 8988 3238
rect 9012 3236 9068 3238
rect 9092 3236 9148 3238
rect 10506 9172 10562 9208
rect 10506 9152 10508 9172
rect 10508 9152 10560 9172
rect 10560 9152 10562 9172
rect 10826 9274 10882 9276
rect 10906 9274 10962 9276
rect 10986 9274 11042 9276
rect 11066 9274 11122 9276
rect 10826 9222 10872 9274
rect 10872 9222 10882 9274
rect 10906 9222 10936 9274
rect 10936 9222 10948 9274
rect 10948 9222 10962 9274
rect 10986 9222 11000 9274
rect 11000 9222 11012 9274
rect 11012 9222 11042 9274
rect 11066 9222 11076 9274
rect 11076 9222 11122 9274
rect 10826 9220 10882 9222
rect 10906 9220 10962 9222
rect 10986 9220 11042 9222
rect 11066 9220 11122 9222
rect 10598 8744 10654 8800
rect 10782 8744 10838 8800
rect 10414 8200 10470 8256
rect 10322 6840 10378 6896
rect 10874 8608 10930 8664
rect 14774 13626 14830 13628
rect 14854 13626 14910 13628
rect 14934 13626 14990 13628
rect 15014 13626 15070 13628
rect 14774 13574 14820 13626
rect 14820 13574 14830 13626
rect 14854 13574 14884 13626
rect 14884 13574 14896 13626
rect 14896 13574 14910 13626
rect 14934 13574 14948 13626
rect 14948 13574 14960 13626
rect 14960 13574 14990 13626
rect 15014 13574 15024 13626
rect 15024 13574 15070 13626
rect 14774 13572 14830 13574
rect 14854 13572 14910 13574
rect 14934 13572 14990 13574
rect 15014 13572 15070 13574
rect 12800 13082 12856 13084
rect 12880 13082 12936 13084
rect 12960 13082 13016 13084
rect 13040 13082 13096 13084
rect 12800 13030 12846 13082
rect 12846 13030 12856 13082
rect 12880 13030 12910 13082
rect 12910 13030 12922 13082
rect 12922 13030 12936 13082
rect 12960 13030 12974 13082
rect 12974 13030 12986 13082
rect 12986 13030 13016 13082
rect 13040 13030 13050 13082
rect 13050 13030 13096 13082
rect 12800 13028 12856 13030
rect 12880 13028 12936 13030
rect 12960 13028 13016 13030
rect 13040 13028 13096 13030
rect 11518 12180 11520 12200
rect 11520 12180 11572 12200
rect 11572 12180 11574 12200
rect 11518 12144 11574 12180
rect 11702 10784 11758 10840
rect 11058 8880 11114 8936
rect 11242 8880 11298 8936
rect 10826 8186 10882 8188
rect 10906 8186 10962 8188
rect 10986 8186 11042 8188
rect 11066 8186 11122 8188
rect 10826 8134 10872 8186
rect 10872 8134 10882 8186
rect 10906 8134 10936 8186
rect 10936 8134 10948 8186
rect 10948 8134 10962 8186
rect 10986 8134 11000 8186
rect 11000 8134 11012 8186
rect 11012 8134 11042 8186
rect 11066 8134 11076 8186
rect 11076 8134 11122 8186
rect 10826 8132 10882 8134
rect 10906 8132 10962 8134
rect 10986 8132 11042 8134
rect 11066 8132 11122 8134
rect 11242 8336 11298 8392
rect 10826 7098 10882 7100
rect 10906 7098 10962 7100
rect 10986 7098 11042 7100
rect 11066 7098 11122 7100
rect 10826 7046 10872 7098
rect 10872 7046 10882 7098
rect 10906 7046 10936 7098
rect 10936 7046 10948 7098
rect 10948 7046 10962 7098
rect 10986 7046 11000 7098
rect 11000 7046 11012 7098
rect 11012 7046 11042 7098
rect 11066 7046 11076 7098
rect 11076 7046 11122 7098
rect 10826 7044 10882 7046
rect 10906 7044 10962 7046
rect 10986 7044 11042 7046
rect 11066 7044 11122 7046
rect 10826 6010 10882 6012
rect 10906 6010 10962 6012
rect 10986 6010 11042 6012
rect 11066 6010 11122 6012
rect 10826 5958 10872 6010
rect 10872 5958 10882 6010
rect 10906 5958 10936 6010
rect 10936 5958 10948 6010
rect 10948 5958 10962 6010
rect 10986 5958 11000 6010
rect 11000 5958 11012 6010
rect 11012 5958 11042 6010
rect 11066 5958 11076 6010
rect 11076 5958 11122 6010
rect 10826 5956 10882 5958
rect 10906 5956 10962 5958
rect 10986 5956 11042 5958
rect 11066 5956 11122 5958
rect 10826 4922 10882 4924
rect 10906 4922 10962 4924
rect 10986 4922 11042 4924
rect 11066 4922 11122 4924
rect 10826 4870 10872 4922
rect 10872 4870 10882 4922
rect 10906 4870 10936 4922
rect 10936 4870 10948 4922
rect 10948 4870 10962 4922
rect 10986 4870 11000 4922
rect 11000 4870 11012 4922
rect 11012 4870 11042 4922
rect 11066 4870 11076 4922
rect 11076 4870 11122 4922
rect 10826 4868 10882 4870
rect 10906 4868 10962 4870
rect 10986 4868 11042 4870
rect 11066 4868 11122 4870
rect 10826 3834 10882 3836
rect 10906 3834 10962 3836
rect 10986 3834 11042 3836
rect 11066 3834 11122 3836
rect 10826 3782 10872 3834
rect 10872 3782 10882 3834
rect 10906 3782 10936 3834
rect 10936 3782 10948 3834
rect 10948 3782 10962 3834
rect 10986 3782 11000 3834
rect 11000 3782 11012 3834
rect 11012 3782 11042 3834
rect 11066 3782 11076 3834
rect 11076 3782 11122 3834
rect 10826 3780 10882 3782
rect 10906 3780 10962 3782
rect 10986 3780 11042 3782
rect 11066 3780 11122 3782
rect 12254 12688 12310 12744
rect 11886 9968 11942 10024
rect 11794 9832 11850 9888
rect 11794 9016 11850 9072
rect 12070 10956 12072 10976
rect 12072 10956 12124 10976
rect 12124 10956 12126 10976
rect 12070 10920 12126 10956
rect 14774 12538 14830 12540
rect 14854 12538 14910 12540
rect 14934 12538 14990 12540
rect 15014 12538 15070 12540
rect 14774 12486 14820 12538
rect 14820 12486 14830 12538
rect 14854 12486 14884 12538
rect 14884 12486 14896 12538
rect 14896 12486 14910 12538
rect 14934 12486 14948 12538
rect 14948 12486 14960 12538
rect 14960 12486 14990 12538
rect 15014 12486 15024 12538
rect 15024 12486 15070 12538
rect 14774 12484 14830 12486
rect 14854 12484 14910 12486
rect 14934 12484 14990 12486
rect 15014 12484 15070 12486
rect 12800 11994 12856 11996
rect 12880 11994 12936 11996
rect 12960 11994 13016 11996
rect 13040 11994 13096 11996
rect 12800 11942 12846 11994
rect 12846 11942 12856 11994
rect 12880 11942 12910 11994
rect 12910 11942 12922 11994
rect 12922 11942 12936 11994
rect 12960 11942 12974 11994
rect 12974 11942 12986 11994
rect 12986 11942 13016 11994
rect 13040 11942 13050 11994
rect 13050 11942 13096 11994
rect 12800 11940 12856 11942
rect 12880 11940 12936 11942
rect 12960 11940 13016 11942
rect 13040 11940 13096 11942
rect 13910 11736 13966 11792
rect 12438 11192 12494 11248
rect 11978 9016 12034 9072
rect 11702 6296 11758 6352
rect 12162 8472 12218 8528
rect 12346 9580 12402 9616
rect 12346 9560 12348 9580
rect 12348 9560 12400 9580
rect 12400 9560 12402 9580
rect 12438 9424 12494 9480
rect 13450 11056 13506 11112
rect 12800 10906 12856 10908
rect 12880 10906 12936 10908
rect 12960 10906 13016 10908
rect 13040 10906 13096 10908
rect 12800 10854 12846 10906
rect 12846 10854 12856 10906
rect 12880 10854 12910 10906
rect 12910 10854 12922 10906
rect 12922 10854 12936 10906
rect 12960 10854 12974 10906
rect 12974 10854 12986 10906
rect 12986 10854 13016 10906
rect 13040 10854 13050 10906
rect 13050 10854 13096 10906
rect 12800 10852 12856 10854
rect 12880 10852 12936 10854
rect 12960 10852 13016 10854
rect 13040 10852 13096 10854
rect 12530 7248 12586 7304
rect 12800 9818 12856 9820
rect 12880 9818 12936 9820
rect 12960 9818 13016 9820
rect 13040 9818 13096 9820
rect 12800 9766 12846 9818
rect 12846 9766 12856 9818
rect 12880 9766 12910 9818
rect 12910 9766 12922 9818
rect 12922 9766 12936 9818
rect 12960 9766 12974 9818
rect 12974 9766 12986 9818
rect 12986 9766 13016 9818
rect 13040 9766 13050 9818
rect 13050 9766 13096 9818
rect 12800 9764 12856 9766
rect 12880 9764 12936 9766
rect 12960 9764 13016 9766
rect 13040 9764 13096 9766
rect 12800 8730 12856 8732
rect 12880 8730 12936 8732
rect 12960 8730 13016 8732
rect 13040 8730 13096 8732
rect 12800 8678 12846 8730
rect 12846 8678 12856 8730
rect 12880 8678 12910 8730
rect 12910 8678 12922 8730
rect 12922 8678 12936 8730
rect 12960 8678 12974 8730
rect 12974 8678 12986 8730
rect 12986 8678 13016 8730
rect 13040 8678 13050 8730
rect 13050 8678 13096 8730
rect 12800 8676 12856 8678
rect 12880 8676 12936 8678
rect 12960 8676 13016 8678
rect 13040 8676 13096 8678
rect 14774 11450 14830 11452
rect 14854 11450 14910 11452
rect 14934 11450 14990 11452
rect 15014 11450 15070 11452
rect 14774 11398 14820 11450
rect 14820 11398 14830 11450
rect 14854 11398 14884 11450
rect 14884 11398 14896 11450
rect 14896 11398 14910 11450
rect 14934 11398 14948 11450
rect 14948 11398 14960 11450
rect 14960 11398 14990 11450
rect 15014 11398 15024 11450
rect 15024 11398 15070 11450
rect 14774 11396 14830 11398
rect 14854 11396 14910 11398
rect 14934 11396 14990 11398
rect 15014 11396 15070 11398
rect 13818 10668 13874 10704
rect 13818 10648 13820 10668
rect 13820 10648 13872 10668
rect 13872 10648 13874 10668
rect 14462 10104 14518 10160
rect 14774 10362 14830 10364
rect 14854 10362 14910 10364
rect 14934 10362 14990 10364
rect 15014 10362 15070 10364
rect 14774 10310 14820 10362
rect 14820 10310 14830 10362
rect 14854 10310 14884 10362
rect 14884 10310 14896 10362
rect 14896 10310 14910 10362
rect 14934 10310 14948 10362
rect 14948 10310 14960 10362
rect 14960 10310 14990 10362
rect 15014 10310 15024 10362
rect 15024 10310 15070 10362
rect 14774 10308 14830 10310
rect 14854 10308 14910 10310
rect 14934 10308 14990 10310
rect 15014 10308 15070 10310
rect 14774 9274 14830 9276
rect 14854 9274 14910 9276
rect 14934 9274 14990 9276
rect 15014 9274 15070 9276
rect 14774 9222 14820 9274
rect 14820 9222 14830 9274
rect 14854 9222 14884 9274
rect 14884 9222 14896 9274
rect 14896 9222 14910 9274
rect 14934 9222 14948 9274
rect 14948 9222 14960 9274
rect 14960 9222 14990 9274
rect 15014 9222 15024 9274
rect 15024 9222 15070 9274
rect 14774 9220 14830 9222
rect 14854 9220 14910 9222
rect 14934 9220 14990 9222
rect 15014 9220 15070 9222
rect 14774 8186 14830 8188
rect 14854 8186 14910 8188
rect 14934 8186 14990 8188
rect 15014 8186 15070 8188
rect 14774 8134 14820 8186
rect 14820 8134 14830 8186
rect 14854 8134 14884 8186
rect 14884 8134 14896 8186
rect 14896 8134 14910 8186
rect 14934 8134 14948 8186
rect 14948 8134 14960 8186
rect 14960 8134 14990 8186
rect 15014 8134 15024 8186
rect 15024 8134 15070 8186
rect 14774 8132 14830 8134
rect 14854 8132 14910 8134
rect 14934 8132 14990 8134
rect 15014 8132 15070 8134
rect 13542 7928 13598 7984
rect 12800 7642 12856 7644
rect 12880 7642 12936 7644
rect 12960 7642 13016 7644
rect 13040 7642 13096 7644
rect 12800 7590 12846 7642
rect 12846 7590 12856 7642
rect 12880 7590 12910 7642
rect 12910 7590 12922 7642
rect 12922 7590 12936 7642
rect 12960 7590 12974 7642
rect 12974 7590 12986 7642
rect 12986 7590 13016 7642
rect 13040 7590 13050 7642
rect 13050 7590 13096 7642
rect 12800 7588 12856 7590
rect 12880 7588 12936 7590
rect 12960 7588 13016 7590
rect 13040 7588 13096 7590
rect 14774 7098 14830 7100
rect 14854 7098 14910 7100
rect 14934 7098 14990 7100
rect 15014 7098 15070 7100
rect 14774 7046 14820 7098
rect 14820 7046 14830 7098
rect 14854 7046 14884 7098
rect 14884 7046 14896 7098
rect 14896 7046 14910 7098
rect 14934 7046 14948 7098
rect 14948 7046 14960 7098
rect 14960 7046 14990 7098
rect 15014 7046 15024 7098
rect 15024 7046 15070 7098
rect 14774 7044 14830 7046
rect 14854 7044 14910 7046
rect 14934 7044 14990 7046
rect 15014 7044 15070 7046
rect 12714 6704 12770 6760
rect 12800 6554 12856 6556
rect 12880 6554 12936 6556
rect 12960 6554 13016 6556
rect 13040 6554 13096 6556
rect 12800 6502 12846 6554
rect 12846 6502 12856 6554
rect 12880 6502 12910 6554
rect 12910 6502 12922 6554
rect 12922 6502 12936 6554
rect 12960 6502 12974 6554
rect 12974 6502 12986 6554
rect 12986 6502 13016 6554
rect 13040 6502 13050 6554
rect 13050 6502 13096 6554
rect 12800 6500 12856 6502
rect 12880 6500 12936 6502
rect 12960 6500 13016 6502
rect 13040 6500 13096 6502
rect 14774 6010 14830 6012
rect 14854 6010 14910 6012
rect 14934 6010 14990 6012
rect 15014 6010 15070 6012
rect 14774 5958 14820 6010
rect 14820 5958 14830 6010
rect 14854 5958 14884 6010
rect 14884 5958 14896 6010
rect 14896 5958 14910 6010
rect 14934 5958 14948 6010
rect 14948 5958 14960 6010
rect 14960 5958 14990 6010
rect 15014 5958 15024 6010
rect 15024 5958 15070 6010
rect 14774 5956 14830 5958
rect 14854 5956 14910 5958
rect 14934 5956 14990 5958
rect 15014 5956 15070 5958
rect 12800 5466 12856 5468
rect 12880 5466 12936 5468
rect 12960 5466 13016 5468
rect 13040 5466 13096 5468
rect 12800 5414 12846 5466
rect 12846 5414 12856 5466
rect 12880 5414 12910 5466
rect 12910 5414 12922 5466
rect 12922 5414 12936 5466
rect 12960 5414 12974 5466
rect 12974 5414 12986 5466
rect 12986 5414 13016 5466
rect 13040 5414 13050 5466
rect 13050 5414 13096 5466
rect 12800 5412 12856 5414
rect 12880 5412 12936 5414
rect 12960 5412 13016 5414
rect 13040 5412 13096 5414
rect 14774 4922 14830 4924
rect 14854 4922 14910 4924
rect 14934 4922 14990 4924
rect 15014 4922 15070 4924
rect 14774 4870 14820 4922
rect 14820 4870 14830 4922
rect 14854 4870 14884 4922
rect 14884 4870 14896 4922
rect 14896 4870 14910 4922
rect 14934 4870 14948 4922
rect 14948 4870 14960 4922
rect 14960 4870 14990 4922
rect 15014 4870 15024 4922
rect 15024 4870 15070 4922
rect 14774 4868 14830 4870
rect 14854 4868 14910 4870
rect 14934 4868 14990 4870
rect 15014 4868 15070 4870
rect 12800 4378 12856 4380
rect 12880 4378 12936 4380
rect 12960 4378 13016 4380
rect 13040 4378 13096 4380
rect 12800 4326 12846 4378
rect 12846 4326 12856 4378
rect 12880 4326 12910 4378
rect 12910 4326 12922 4378
rect 12922 4326 12936 4378
rect 12960 4326 12974 4378
rect 12974 4326 12986 4378
rect 12986 4326 13016 4378
rect 13040 4326 13050 4378
rect 13050 4326 13096 4378
rect 12800 4324 12856 4326
rect 12880 4324 12936 4326
rect 12960 4324 13016 4326
rect 13040 4324 13096 4326
rect 14774 3834 14830 3836
rect 14854 3834 14910 3836
rect 14934 3834 14990 3836
rect 15014 3834 15070 3836
rect 14774 3782 14820 3834
rect 14820 3782 14830 3834
rect 14854 3782 14884 3834
rect 14884 3782 14896 3834
rect 14896 3782 14910 3834
rect 14934 3782 14948 3834
rect 14948 3782 14960 3834
rect 14960 3782 14990 3834
rect 15014 3782 15024 3834
rect 15024 3782 15070 3834
rect 14774 3780 14830 3782
rect 14854 3780 14910 3782
rect 14934 3780 14990 3782
rect 15014 3780 15070 3782
rect 12800 3290 12856 3292
rect 12880 3290 12936 3292
rect 12960 3290 13016 3292
rect 13040 3290 13096 3292
rect 12800 3238 12846 3290
rect 12846 3238 12856 3290
rect 12880 3238 12910 3290
rect 12910 3238 12922 3290
rect 12922 3238 12936 3290
rect 12960 3238 12974 3290
rect 12974 3238 12986 3290
rect 12986 3238 13016 3290
rect 13040 3238 13050 3290
rect 13050 3238 13096 3290
rect 12800 3236 12856 3238
rect 12880 3236 12936 3238
rect 12960 3236 13016 3238
rect 13040 3236 13096 3238
rect 6878 2746 6934 2748
rect 6958 2746 7014 2748
rect 7038 2746 7094 2748
rect 7118 2746 7174 2748
rect 6878 2694 6924 2746
rect 6924 2694 6934 2746
rect 6958 2694 6988 2746
rect 6988 2694 7000 2746
rect 7000 2694 7014 2746
rect 7038 2694 7052 2746
rect 7052 2694 7064 2746
rect 7064 2694 7094 2746
rect 7118 2694 7128 2746
rect 7128 2694 7174 2746
rect 6878 2692 6934 2694
rect 6958 2692 7014 2694
rect 7038 2692 7094 2694
rect 7118 2692 7174 2694
rect 10826 2746 10882 2748
rect 10906 2746 10962 2748
rect 10986 2746 11042 2748
rect 11066 2746 11122 2748
rect 10826 2694 10872 2746
rect 10872 2694 10882 2746
rect 10906 2694 10936 2746
rect 10936 2694 10948 2746
rect 10948 2694 10962 2746
rect 10986 2694 11000 2746
rect 11000 2694 11012 2746
rect 11012 2694 11042 2746
rect 11066 2694 11076 2746
rect 11076 2694 11122 2746
rect 10826 2692 10882 2694
rect 10906 2692 10962 2694
rect 10986 2692 11042 2694
rect 11066 2692 11122 2694
rect 14774 2746 14830 2748
rect 14854 2746 14910 2748
rect 14934 2746 14990 2748
rect 15014 2746 15070 2748
rect 14774 2694 14820 2746
rect 14820 2694 14830 2746
rect 14854 2694 14884 2746
rect 14884 2694 14896 2746
rect 14896 2694 14910 2746
rect 14934 2694 14948 2746
rect 14948 2694 14960 2746
rect 14960 2694 14990 2746
rect 15014 2694 15024 2746
rect 15024 2694 15070 2746
rect 14774 2692 14830 2694
rect 14854 2692 14910 2694
rect 14934 2692 14990 2694
rect 15014 2692 15070 2694
rect 4904 2202 4960 2204
rect 4984 2202 5040 2204
rect 5064 2202 5120 2204
rect 5144 2202 5200 2204
rect 4904 2150 4950 2202
rect 4950 2150 4960 2202
rect 4984 2150 5014 2202
rect 5014 2150 5026 2202
rect 5026 2150 5040 2202
rect 5064 2150 5078 2202
rect 5078 2150 5090 2202
rect 5090 2150 5120 2202
rect 5144 2150 5154 2202
rect 5154 2150 5200 2202
rect 4904 2148 4960 2150
rect 4984 2148 5040 2150
rect 5064 2148 5120 2150
rect 5144 2148 5200 2150
rect 8852 2202 8908 2204
rect 8932 2202 8988 2204
rect 9012 2202 9068 2204
rect 9092 2202 9148 2204
rect 8852 2150 8898 2202
rect 8898 2150 8908 2202
rect 8932 2150 8962 2202
rect 8962 2150 8974 2202
rect 8974 2150 8988 2202
rect 9012 2150 9026 2202
rect 9026 2150 9038 2202
rect 9038 2150 9068 2202
rect 9092 2150 9102 2202
rect 9102 2150 9148 2202
rect 8852 2148 8908 2150
rect 8932 2148 8988 2150
rect 9012 2148 9068 2150
rect 9092 2148 9148 2150
rect 12800 2202 12856 2204
rect 12880 2202 12936 2204
rect 12960 2202 13016 2204
rect 13040 2202 13096 2204
rect 12800 2150 12846 2202
rect 12846 2150 12856 2202
rect 12880 2150 12910 2202
rect 12910 2150 12922 2202
rect 12922 2150 12936 2202
rect 12960 2150 12974 2202
rect 12974 2150 12986 2202
rect 12986 2150 13016 2202
rect 13040 2150 13050 2202
rect 13050 2150 13096 2202
rect 12800 2148 12856 2150
rect 12880 2148 12936 2150
rect 12960 2148 13016 2150
rect 13040 2148 13096 2150
rect 2930 1658 2986 1660
rect 3010 1658 3066 1660
rect 3090 1658 3146 1660
rect 3170 1658 3226 1660
rect 2930 1606 2976 1658
rect 2976 1606 2986 1658
rect 3010 1606 3040 1658
rect 3040 1606 3052 1658
rect 3052 1606 3066 1658
rect 3090 1606 3104 1658
rect 3104 1606 3116 1658
rect 3116 1606 3146 1658
rect 3170 1606 3180 1658
rect 3180 1606 3226 1658
rect 2930 1604 2986 1606
rect 3010 1604 3066 1606
rect 3090 1604 3146 1606
rect 3170 1604 3226 1606
rect 6878 1658 6934 1660
rect 6958 1658 7014 1660
rect 7038 1658 7094 1660
rect 7118 1658 7174 1660
rect 6878 1606 6924 1658
rect 6924 1606 6934 1658
rect 6958 1606 6988 1658
rect 6988 1606 7000 1658
rect 7000 1606 7014 1658
rect 7038 1606 7052 1658
rect 7052 1606 7064 1658
rect 7064 1606 7094 1658
rect 7118 1606 7128 1658
rect 7128 1606 7174 1658
rect 6878 1604 6934 1606
rect 6958 1604 7014 1606
rect 7038 1604 7094 1606
rect 7118 1604 7174 1606
rect 10826 1658 10882 1660
rect 10906 1658 10962 1660
rect 10986 1658 11042 1660
rect 11066 1658 11122 1660
rect 10826 1606 10872 1658
rect 10872 1606 10882 1658
rect 10906 1606 10936 1658
rect 10936 1606 10948 1658
rect 10948 1606 10962 1658
rect 10986 1606 11000 1658
rect 11000 1606 11012 1658
rect 11012 1606 11042 1658
rect 11066 1606 11076 1658
rect 11076 1606 11122 1658
rect 10826 1604 10882 1606
rect 10906 1604 10962 1606
rect 10986 1604 11042 1606
rect 11066 1604 11122 1606
rect 14774 1658 14830 1660
rect 14854 1658 14910 1660
rect 14934 1658 14990 1660
rect 15014 1658 15070 1660
rect 14774 1606 14820 1658
rect 14820 1606 14830 1658
rect 14854 1606 14884 1658
rect 14884 1606 14896 1658
rect 14896 1606 14910 1658
rect 14934 1606 14948 1658
rect 14948 1606 14960 1658
rect 14960 1606 14990 1658
rect 15014 1606 15024 1658
rect 15024 1606 15070 1658
rect 14774 1604 14830 1606
rect 14854 1604 14910 1606
rect 14934 1604 14990 1606
rect 15014 1604 15070 1606
rect 4904 1114 4960 1116
rect 4984 1114 5040 1116
rect 5064 1114 5120 1116
rect 5144 1114 5200 1116
rect 4904 1062 4950 1114
rect 4950 1062 4960 1114
rect 4984 1062 5014 1114
rect 5014 1062 5026 1114
rect 5026 1062 5040 1114
rect 5064 1062 5078 1114
rect 5078 1062 5090 1114
rect 5090 1062 5120 1114
rect 5144 1062 5154 1114
rect 5154 1062 5200 1114
rect 4904 1060 4960 1062
rect 4984 1060 5040 1062
rect 5064 1060 5120 1062
rect 5144 1060 5200 1062
rect 8852 1114 8908 1116
rect 8932 1114 8988 1116
rect 9012 1114 9068 1116
rect 9092 1114 9148 1116
rect 8852 1062 8898 1114
rect 8898 1062 8908 1114
rect 8932 1062 8962 1114
rect 8962 1062 8974 1114
rect 8974 1062 8988 1114
rect 9012 1062 9026 1114
rect 9026 1062 9038 1114
rect 9038 1062 9068 1114
rect 9092 1062 9102 1114
rect 9102 1062 9148 1114
rect 8852 1060 8908 1062
rect 8932 1060 8988 1062
rect 9012 1060 9068 1062
rect 9092 1060 9148 1062
rect 12800 1114 12856 1116
rect 12880 1114 12936 1116
rect 12960 1114 13016 1116
rect 13040 1114 13096 1116
rect 12800 1062 12846 1114
rect 12846 1062 12856 1114
rect 12880 1062 12910 1114
rect 12910 1062 12922 1114
rect 12922 1062 12936 1114
rect 12960 1062 12974 1114
rect 12974 1062 12986 1114
rect 12986 1062 13016 1114
rect 13040 1062 13050 1114
rect 13050 1062 13096 1114
rect 12800 1060 12856 1062
rect 12880 1060 12936 1062
rect 12960 1060 13016 1062
rect 13040 1060 13096 1062
rect 1398 720 1454 776
<< metal3 >>
rect 0 23218 400 23248
rect 2773 23218 2839 23221
rect 0 23216 2839 23218
rect 0 23160 2778 23216
rect 2834 23160 2839 23216
rect 0 23158 2839 23160
rect 0 23128 400 23158
rect 2773 23155 2839 23158
rect 4894 22880 5210 22881
rect 4894 22816 4900 22880
rect 4964 22816 4980 22880
rect 5044 22816 5060 22880
rect 5124 22816 5140 22880
rect 5204 22816 5210 22880
rect 4894 22815 5210 22816
rect 8842 22880 9158 22881
rect 8842 22816 8848 22880
rect 8912 22816 8928 22880
rect 8992 22816 9008 22880
rect 9072 22816 9088 22880
rect 9152 22816 9158 22880
rect 8842 22815 9158 22816
rect 12790 22880 13106 22881
rect 12790 22816 12796 22880
rect 12860 22816 12876 22880
rect 12940 22816 12956 22880
rect 13020 22816 13036 22880
rect 13100 22816 13106 22880
rect 12790 22815 13106 22816
rect 2920 22336 3236 22337
rect 2920 22272 2926 22336
rect 2990 22272 3006 22336
rect 3070 22272 3086 22336
rect 3150 22272 3166 22336
rect 3230 22272 3236 22336
rect 2920 22271 3236 22272
rect 6868 22336 7184 22337
rect 6868 22272 6874 22336
rect 6938 22272 6954 22336
rect 7018 22272 7034 22336
rect 7098 22272 7114 22336
rect 7178 22272 7184 22336
rect 6868 22271 7184 22272
rect 10816 22336 11132 22337
rect 10816 22272 10822 22336
rect 10886 22272 10902 22336
rect 10966 22272 10982 22336
rect 11046 22272 11062 22336
rect 11126 22272 11132 22336
rect 10816 22271 11132 22272
rect 14764 22336 15080 22337
rect 14764 22272 14770 22336
rect 14834 22272 14850 22336
rect 14914 22272 14930 22336
rect 14994 22272 15010 22336
rect 15074 22272 15080 22336
rect 14764 22271 15080 22272
rect 4894 21792 5210 21793
rect 0 21722 400 21752
rect 4894 21728 4900 21792
rect 4964 21728 4980 21792
rect 5044 21728 5060 21792
rect 5124 21728 5140 21792
rect 5204 21728 5210 21792
rect 4894 21727 5210 21728
rect 8842 21792 9158 21793
rect 8842 21728 8848 21792
rect 8912 21728 8928 21792
rect 8992 21728 9008 21792
rect 9072 21728 9088 21792
rect 9152 21728 9158 21792
rect 8842 21727 9158 21728
rect 12790 21792 13106 21793
rect 12790 21728 12796 21792
rect 12860 21728 12876 21792
rect 12940 21728 12956 21792
rect 13020 21728 13036 21792
rect 13100 21728 13106 21792
rect 12790 21727 13106 21728
rect 1485 21722 1551 21725
rect 0 21720 1551 21722
rect 0 21664 1490 21720
rect 1546 21664 1551 21720
rect 0 21662 1551 21664
rect 0 21632 400 21662
rect 1485 21659 1551 21662
rect 2920 21248 3236 21249
rect 2920 21184 2926 21248
rect 2990 21184 3006 21248
rect 3070 21184 3086 21248
rect 3150 21184 3166 21248
rect 3230 21184 3236 21248
rect 2920 21183 3236 21184
rect 6868 21248 7184 21249
rect 6868 21184 6874 21248
rect 6938 21184 6954 21248
rect 7018 21184 7034 21248
rect 7098 21184 7114 21248
rect 7178 21184 7184 21248
rect 6868 21183 7184 21184
rect 10816 21248 11132 21249
rect 10816 21184 10822 21248
rect 10886 21184 10902 21248
rect 10966 21184 10982 21248
rect 11046 21184 11062 21248
rect 11126 21184 11132 21248
rect 10816 21183 11132 21184
rect 14764 21248 15080 21249
rect 14764 21184 14770 21248
rect 14834 21184 14850 21248
rect 14914 21184 14930 21248
rect 14994 21184 15010 21248
rect 15074 21184 15080 21248
rect 14764 21183 15080 21184
rect 4894 20704 5210 20705
rect 4894 20640 4900 20704
rect 4964 20640 4980 20704
rect 5044 20640 5060 20704
rect 5124 20640 5140 20704
rect 5204 20640 5210 20704
rect 4894 20639 5210 20640
rect 8842 20704 9158 20705
rect 8842 20640 8848 20704
rect 8912 20640 8928 20704
rect 8992 20640 9008 20704
rect 9072 20640 9088 20704
rect 9152 20640 9158 20704
rect 8842 20639 9158 20640
rect 12790 20704 13106 20705
rect 12790 20640 12796 20704
rect 12860 20640 12876 20704
rect 12940 20640 12956 20704
rect 13020 20640 13036 20704
rect 13100 20640 13106 20704
rect 12790 20639 13106 20640
rect 0 20226 400 20256
rect 0 20166 2790 20226
rect 0 20136 400 20166
rect 2730 19954 2790 20166
rect 2920 20160 3236 20161
rect 2920 20096 2926 20160
rect 2990 20096 3006 20160
rect 3070 20096 3086 20160
rect 3150 20096 3166 20160
rect 3230 20096 3236 20160
rect 2920 20095 3236 20096
rect 6868 20160 7184 20161
rect 6868 20096 6874 20160
rect 6938 20096 6954 20160
rect 7018 20096 7034 20160
rect 7098 20096 7114 20160
rect 7178 20096 7184 20160
rect 6868 20095 7184 20096
rect 10816 20160 11132 20161
rect 10816 20096 10822 20160
rect 10886 20096 10902 20160
rect 10966 20096 10982 20160
rect 11046 20096 11062 20160
rect 11126 20096 11132 20160
rect 10816 20095 11132 20096
rect 14764 20160 15080 20161
rect 14764 20096 14770 20160
rect 14834 20096 14850 20160
rect 14914 20096 14930 20160
rect 14994 20096 15010 20160
rect 15074 20096 15080 20160
rect 14764 20095 15080 20096
rect 3325 19954 3391 19957
rect 2730 19952 3391 19954
rect 2730 19896 3330 19952
rect 3386 19896 3391 19952
rect 2730 19894 3391 19896
rect 3325 19891 3391 19894
rect 4894 19616 5210 19617
rect 4894 19552 4900 19616
rect 4964 19552 4980 19616
rect 5044 19552 5060 19616
rect 5124 19552 5140 19616
rect 5204 19552 5210 19616
rect 4894 19551 5210 19552
rect 8842 19616 9158 19617
rect 8842 19552 8848 19616
rect 8912 19552 8928 19616
rect 8992 19552 9008 19616
rect 9072 19552 9088 19616
rect 9152 19552 9158 19616
rect 8842 19551 9158 19552
rect 12790 19616 13106 19617
rect 12790 19552 12796 19616
rect 12860 19552 12876 19616
rect 12940 19552 12956 19616
rect 13020 19552 13036 19616
rect 13100 19552 13106 19616
rect 12790 19551 13106 19552
rect 2920 19072 3236 19073
rect 2920 19008 2926 19072
rect 2990 19008 3006 19072
rect 3070 19008 3086 19072
rect 3150 19008 3166 19072
rect 3230 19008 3236 19072
rect 2920 19007 3236 19008
rect 6868 19072 7184 19073
rect 6868 19008 6874 19072
rect 6938 19008 6954 19072
rect 7018 19008 7034 19072
rect 7098 19008 7114 19072
rect 7178 19008 7184 19072
rect 6868 19007 7184 19008
rect 10816 19072 11132 19073
rect 10816 19008 10822 19072
rect 10886 19008 10902 19072
rect 10966 19008 10982 19072
rect 11046 19008 11062 19072
rect 11126 19008 11132 19072
rect 10816 19007 11132 19008
rect 14764 19072 15080 19073
rect 14764 19008 14770 19072
rect 14834 19008 14850 19072
rect 14914 19008 14930 19072
rect 14994 19008 15010 19072
rect 15074 19008 15080 19072
rect 14764 19007 15080 19008
rect 0 18730 400 18760
rect 2773 18730 2839 18733
rect 0 18728 2839 18730
rect 0 18672 2778 18728
rect 2834 18672 2839 18728
rect 0 18670 2839 18672
rect 0 18640 400 18670
rect 2773 18667 2839 18670
rect 4894 18528 5210 18529
rect 4894 18464 4900 18528
rect 4964 18464 4980 18528
rect 5044 18464 5060 18528
rect 5124 18464 5140 18528
rect 5204 18464 5210 18528
rect 4894 18463 5210 18464
rect 8842 18528 9158 18529
rect 8842 18464 8848 18528
rect 8912 18464 8928 18528
rect 8992 18464 9008 18528
rect 9072 18464 9088 18528
rect 9152 18464 9158 18528
rect 8842 18463 9158 18464
rect 12790 18528 13106 18529
rect 12790 18464 12796 18528
rect 12860 18464 12876 18528
rect 12940 18464 12956 18528
rect 13020 18464 13036 18528
rect 13100 18464 13106 18528
rect 12790 18463 13106 18464
rect 2920 17984 3236 17985
rect 2920 17920 2926 17984
rect 2990 17920 3006 17984
rect 3070 17920 3086 17984
rect 3150 17920 3166 17984
rect 3230 17920 3236 17984
rect 2920 17919 3236 17920
rect 6868 17984 7184 17985
rect 6868 17920 6874 17984
rect 6938 17920 6954 17984
rect 7018 17920 7034 17984
rect 7098 17920 7114 17984
rect 7178 17920 7184 17984
rect 6868 17919 7184 17920
rect 10816 17984 11132 17985
rect 10816 17920 10822 17984
rect 10886 17920 10902 17984
rect 10966 17920 10982 17984
rect 11046 17920 11062 17984
rect 11126 17920 11132 17984
rect 10816 17919 11132 17920
rect 14764 17984 15080 17985
rect 14764 17920 14770 17984
rect 14834 17920 14850 17984
rect 14914 17920 14930 17984
rect 14994 17920 15010 17984
rect 15074 17920 15080 17984
rect 14764 17919 15080 17920
rect 4894 17440 5210 17441
rect 4894 17376 4900 17440
rect 4964 17376 4980 17440
rect 5044 17376 5060 17440
rect 5124 17376 5140 17440
rect 5204 17376 5210 17440
rect 4894 17375 5210 17376
rect 8842 17440 9158 17441
rect 8842 17376 8848 17440
rect 8912 17376 8928 17440
rect 8992 17376 9008 17440
rect 9072 17376 9088 17440
rect 9152 17376 9158 17440
rect 8842 17375 9158 17376
rect 12790 17440 13106 17441
rect 12790 17376 12796 17440
rect 12860 17376 12876 17440
rect 12940 17376 12956 17440
rect 13020 17376 13036 17440
rect 13100 17376 13106 17440
rect 12790 17375 13106 17376
rect 0 17234 400 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 400 17174
rect 1485 17171 1551 17174
rect 2920 16896 3236 16897
rect 2920 16832 2926 16896
rect 2990 16832 3006 16896
rect 3070 16832 3086 16896
rect 3150 16832 3166 16896
rect 3230 16832 3236 16896
rect 2920 16831 3236 16832
rect 6868 16896 7184 16897
rect 6868 16832 6874 16896
rect 6938 16832 6954 16896
rect 7018 16832 7034 16896
rect 7098 16832 7114 16896
rect 7178 16832 7184 16896
rect 6868 16831 7184 16832
rect 10816 16896 11132 16897
rect 10816 16832 10822 16896
rect 10886 16832 10902 16896
rect 10966 16832 10982 16896
rect 11046 16832 11062 16896
rect 11126 16832 11132 16896
rect 10816 16831 11132 16832
rect 14764 16896 15080 16897
rect 14764 16832 14770 16896
rect 14834 16832 14850 16896
rect 14914 16832 14930 16896
rect 14994 16832 15010 16896
rect 15074 16832 15080 16896
rect 14764 16831 15080 16832
rect 4894 16352 5210 16353
rect 4894 16288 4900 16352
rect 4964 16288 4980 16352
rect 5044 16288 5060 16352
rect 5124 16288 5140 16352
rect 5204 16288 5210 16352
rect 4894 16287 5210 16288
rect 8842 16352 9158 16353
rect 8842 16288 8848 16352
rect 8912 16288 8928 16352
rect 8992 16288 9008 16352
rect 9072 16288 9088 16352
rect 9152 16288 9158 16352
rect 8842 16287 9158 16288
rect 12790 16352 13106 16353
rect 12790 16288 12796 16352
rect 12860 16288 12876 16352
rect 12940 16288 12956 16352
rect 13020 16288 13036 16352
rect 13100 16288 13106 16352
rect 12790 16287 13106 16288
rect 2920 15808 3236 15809
rect 0 15738 400 15768
rect 2920 15744 2926 15808
rect 2990 15744 3006 15808
rect 3070 15744 3086 15808
rect 3150 15744 3166 15808
rect 3230 15744 3236 15808
rect 2920 15743 3236 15744
rect 6868 15808 7184 15809
rect 6868 15744 6874 15808
rect 6938 15744 6954 15808
rect 7018 15744 7034 15808
rect 7098 15744 7114 15808
rect 7178 15744 7184 15808
rect 6868 15743 7184 15744
rect 10816 15808 11132 15809
rect 10816 15744 10822 15808
rect 10886 15744 10902 15808
rect 10966 15744 10982 15808
rect 11046 15744 11062 15808
rect 11126 15744 11132 15808
rect 10816 15743 11132 15744
rect 14764 15808 15080 15809
rect 14764 15744 14770 15808
rect 14834 15744 14850 15808
rect 14914 15744 14930 15808
rect 14994 15744 15010 15808
rect 15074 15744 15080 15808
rect 14764 15743 15080 15744
rect 2773 15738 2839 15741
rect 0 15736 2839 15738
rect 0 15680 2778 15736
rect 2834 15680 2839 15736
rect 0 15678 2839 15680
rect 0 15648 400 15678
rect 2773 15675 2839 15678
rect 4337 15602 4403 15605
rect 5717 15602 5783 15605
rect 4337 15600 5783 15602
rect 4337 15544 4342 15600
rect 4398 15544 5722 15600
rect 5778 15544 5783 15600
rect 4337 15542 5783 15544
rect 4337 15539 4403 15542
rect 5717 15539 5783 15542
rect 4705 15466 4771 15469
rect 5390 15466 5396 15468
rect 4705 15464 5396 15466
rect 4705 15408 4710 15464
rect 4766 15408 5396 15464
rect 4705 15406 5396 15408
rect 4705 15403 4771 15406
rect 5390 15404 5396 15406
rect 5460 15404 5466 15468
rect 5809 15466 5875 15469
rect 6494 15466 6500 15468
rect 5809 15464 6500 15466
rect 5809 15408 5814 15464
rect 5870 15408 6500 15464
rect 5809 15406 6500 15408
rect 5809 15403 5875 15406
rect 6494 15404 6500 15406
rect 6564 15404 6570 15468
rect 4894 15264 5210 15265
rect 4894 15200 4900 15264
rect 4964 15200 4980 15264
rect 5044 15200 5060 15264
rect 5124 15200 5140 15264
rect 5204 15200 5210 15264
rect 4894 15199 5210 15200
rect 8842 15264 9158 15265
rect 8842 15200 8848 15264
rect 8912 15200 8928 15264
rect 8992 15200 9008 15264
rect 9072 15200 9088 15264
rect 9152 15200 9158 15264
rect 8842 15199 9158 15200
rect 12790 15264 13106 15265
rect 12790 15200 12796 15264
rect 12860 15200 12876 15264
rect 12940 15200 12956 15264
rect 13020 15200 13036 15264
rect 13100 15200 13106 15264
rect 12790 15199 13106 15200
rect 3417 15058 3483 15061
rect 7649 15058 7715 15061
rect 3417 15056 7715 15058
rect 3417 15000 3422 15056
rect 3478 15000 7654 15056
rect 7710 15000 7715 15056
rect 3417 14998 7715 15000
rect 3417 14995 3483 14998
rect 7649 14995 7715 14998
rect 2037 14922 2103 14925
rect 6361 14922 6427 14925
rect 2037 14920 6427 14922
rect 2037 14864 2042 14920
rect 2098 14864 6366 14920
rect 6422 14864 6427 14920
rect 2037 14862 6427 14864
rect 2037 14859 2103 14862
rect 6361 14859 6427 14862
rect 7097 14922 7163 14925
rect 7414 14922 7420 14924
rect 7097 14920 7420 14922
rect 7097 14864 7102 14920
rect 7158 14864 7420 14920
rect 7097 14862 7420 14864
rect 7097 14859 7163 14862
rect 7414 14860 7420 14862
rect 7484 14860 7490 14924
rect 2920 14720 3236 14721
rect 2920 14656 2926 14720
rect 2990 14656 3006 14720
rect 3070 14656 3086 14720
rect 3150 14656 3166 14720
rect 3230 14656 3236 14720
rect 2920 14655 3236 14656
rect 6868 14720 7184 14721
rect 6868 14656 6874 14720
rect 6938 14656 6954 14720
rect 7018 14656 7034 14720
rect 7098 14656 7114 14720
rect 7178 14656 7184 14720
rect 6868 14655 7184 14656
rect 10816 14720 11132 14721
rect 10816 14656 10822 14720
rect 10886 14656 10902 14720
rect 10966 14656 10982 14720
rect 11046 14656 11062 14720
rect 11126 14656 11132 14720
rect 10816 14655 11132 14656
rect 14764 14720 15080 14721
rect 14764 14656 14770 14720
rect 14834 14656 14850 14720
rect 14914 14656 14930 14720
rect 14994 14656 15010 14720
rect 15074 14656 15080 14720
rect 14764 14655 15080 14656
rect 3918 14316 3924 14380
rect 3988 14378 3994 14380
rect 5993 14378 6059 14381
rect 10593 14378 10659 14381
rect 3988 14376 10659 14378
rect 3988 14320 5998 14376
rect 6054 14320 10598 14376
rect 10654 14320 10659 14376
rect 3988 14318 10659 14320
rect 3988 14316 3994 14318
rect 5993 14315 6059 14318
rect 10593 14315 10659 14318
rect 0 14242 400 14272
rect 3325 14242 3391 14245
rect 0 14240 3391 14242
rect 0 14184 3330 14240
rect 3386 14184 3391 14240
rect 0 14182 3391 14184
rect 0 14152 400 14182
rect 3325 14179 3391 14182
rect 4894 14176 5210 14177
rect 4894 14112 4900 14176
rect 4964 14112 4980 14176
rect 5044 14112 5060 14176
rect 5124 14112 5140 14176
rect 5204 14112 5210 14176
rect 4894 14111 5210 14112
rect 8842 14176 9158 14177
rect 8842 14112 8848 14176
rect 8912 14112 8928 14176
rect 8992 14112 9008 14176
rect 9072 14112 9088 14176
rect 9152 14112 9158 14176
rect 8842 14111 9158 14112
rect 12790 14176 13106 14177
rect 12790 14112 12796 14176
rect 12860 14112 12876 14176
rect 12940 14112 12956 14176
rect 13020 14112 13036 14176
rect 13100 14112 13106 14176
rect 12790 14111 13106 14112
rect 5441 14106 5507 14109
rect 7557 14106 7623 14109
rect 5441 14104 7623 14106
rect 5441 14048 5446 14104
rect 5502 14048 7562 14104
rect 7618 14048 7623 14104
rect 5441 14046 7623 14048
rect 5441 14043 5507 14046
rect 7557 14043 7623 14046
rect 5717 13970 5783 13973
rect 10317 13970 10383 13973
rect 5717 13968 10383 13970
rect 5717 13912 5722 13968
rect 5778 13912 10322 13968
rect 10378 13912 10383 13968
rect 5717 13910 10383 13912
rect 5717 13907 5783 13910
rect 10317 13907 10383 13910
rect 2920 13632 3236 13633
rect 2920 13568 2926 13632
rect 2990 13568 3006 13632
rect 3070 13568 3086 13632
rect 3150 13568 3166 13632
rect 3230 13568 3236 13632
rect 2920 13567 3236 13568
rect 6868 13632 7184 13633
rect 6868 13568 6874 13632
rect 6938 13568 6954 13632
rect 7018 13568 7034 13632
rect 7098 13568 7114 13632
rect 7178 13568 7184 13632
rect 6868 13567 7184 13568
rect 10816 13632 11132 13633
rect 10816 13568 10822 13632
rect 10886 13568 10902 13632
rect 10966 13568 10982 13632
rect 11046 13568 11062 13632
rect 11126 13568 11132 13632
rect 10816 13567 11132 13568
rect 14764 13632 15080 13633
rect 14764 13568 14770 13632
rect 14834 13568 14850 13632
rect 14914 13568 14930 13632
rect 14994 13568 15010 13632
rect 15074 13568 15080 13632
rect 14764 13567 15080 13568
rect 3877 13562 3943 13565
rect 3877 13560 3986 13562
rect 3877 13504 3882 13560
rect 3938 13504 3986 13560
rect 3877 13499 3986 13504
rect 2681 13426 2747 13429
rect 3926 13426 3986 13499
rect 6729 13426 6795 13429
rect 2681 13424 6795 13426
rect 2681 13368 2686 13424
rect 2742 13368 6734 13424
rect 6790 13368 6795 13424
rect 2681 13366 6795 13368
rect 2681 13363 2747 13366
rect 6729 13363 6795 13366
rect 8017 13426 8083 13429
rect 8702 13426 8708 13428
rect 8017 13424 8708 13426
rect 8017 13368 8022 13424
rect 8078 13368 8708 13424
rect 8017 13366 8708 13368
rect 8017 13363 8083 13366
rect 8702 13364 8708 13366
rect 8772 13364 8778 13428
rect 2773 13290 2839 13293
rect 8661 13290 8727 13293
rect 2773 13288 8727 13290
rect 2773 13232 2778 13288
rect 2834 13232 8666 13288
rect 8722 13232 8727 13288
rect 2773 13230 8727 13232
rect 2773 13227 2839 13230
rect 8661 13227 8727 13230
rect 4894 13088 5210 13089
rect 4894 13024 4900 13088
rect 4964 13024 4980 13088
rect 5044 13024 5060 13088
rect 5124 13024 5140 13088
rect 5204 13024 5210 13088
rect 4894 13023 5210 13024
rect 8842 13088 9158 13089
rect 8842 13024 8848 13088
rect 8912 13024 8928 13088
rect 8992 13024 9008 13088
rect 9072 13024 9088 13088
rect 9152 13024 9158 13088
rect 8842 13023 9158 13024
rect 12790 13088 13106 13089
rect 12790 13024 12796 13088
rect 12860 13024 12876 13088
rect 12940 13024 12956 13088
rect 13020 13024 13036 13088
rect 13100 13024 13106 13088
rect 12790 13023 13106 13024
rect 2957 12882 3023 12885
rect 4705 12882 4771 12885
rect 8109 12882 8175 12885
rect 10133 12882 10199 12885
rect 2957 12880 3802 12882
rect 2957 12824 2962 12880
rect 3018 12824 3802 12880
rect 2957 12822 3802 12824
rect 2957 12819 3023 12822
rect 0 12746 400 12776
rect 3509 12746 3575 12749
rect 0 12744 3575 12746
rect 0 12688 3514 12744
rect 3570 12688 3575 12744
rect 0 12686 3575 12688
rect 3742 12746 3802 12822
rect 4705 12880 10199 12882
rect 4705 12824 4710 12880
rect 4766 12824 8114 12880
rect 8170 12824 10138 12880
rect 10194 12824 10199 12880
rect 4705 12822 10199 12824
rect 4705 12819 4771 12822
rect 8109 12819 8175 12822
rect 10133 12819 10199 12822
rect 5533 12746 5599 12749
rect 3742 12744 5599 12746
rect 3742 12688 5538 12744
rect 5594 12688 5599 12744
rect 3742 12686 5599 12688
rect 0 12656 400 12686
rect 3509 12683 3575 12686
rect 5533 12683 5599 12686
rect 9029 12746 9095 12749
rect 12249 12746 12315 12749
rect 9029 12744 12315 12746
rect 9029 12688 9034 12744
rect 9090 12688 12254 12744
rect 12310 12688 12315 12744
rect 9029 12686 12315 12688
rect 9029 12683 9095 12686
rect 12249 12683 12315 12686
rect 3417 12610 3483 12613
rect 4981 12610 5047 12613
rect 3417 12608 5047 12610
rect 3417 12552 3422 12608
rect 3478 12552 4986 12608
rect 5042 12552 5047 12608
rect 3417 12550 5047 12552
rect 3417 12547 3483 12550
rect 4981 12547 5047 12550
rect 8017 12610 8083 12613
rect 8017 12608 10012 12610
rect 8017 12552 8022 12608
rect 8078 12552 10012 12608
rect 8017 12550 10012 12552
rect 8017 12547 8083 12550
rect 2920 12544 3236 12545
rect 2920 12480 2926 12544
rect 2990 12480 3006 12544
rect 3070 12480 3086 12544
rect 3150 12480 3166 12544
rect 3230 12480 3236 12544
rect 2920 12479 3236 12480
rect 6868 12544 7184 12545
rect 6868 12480 6874 12544
rect 6938 12480 6954 12544
rect 7018 12480 7034 12544
rect 7098 12480 7114 12544
rect 7178 12480 7184 12544
rect 6868 12479 7184 12480
rect 8845 12474 8911 12477
rect 9489 12476 9555 12477
rect 9254 12474 9260 12476
rect 8845 12472 9260 12474
rect 8845 12416 8850 12472
rect 8906 12416 9260 12472
rect 8845 12414 9260 12416
rect 8845 12411 8911 12414
rect 9254 12412 9260 12414
rect 9324 12412 9330 12476
rect 9438 12474 9444 12476
rect 9398 12414 9444 12474
rect 9508 12472 9555 12476
rect 9550 12416 9555 12472
rect 9438 12412 9444 12414
rect 9508 12412 9555 12416
rect 9489 12411 9555 12412
rect 2497 12338 2563 12341
rect 6729 12338 6795 12341
rect 9121 12338 9187 12341
rect 2497 12336 9187 12338
rect 2497 12280 2502 12336
rect 2558 12280 6734 12336
rect 6790 12280 9126 12336
rect 9182 12280 9187 12336
rect 2497 12278 9187 12280
rect 2497 12275 2563 12278
rect 6729 12275 6795 12278
rect 9121 12275 9187 12278
rect 9673 12338 9739 12341
rect 9806 12338 9812 12340
rect 9673 12336 9812 12338
rect 9673 12280 9678 12336
rect 9734 12280 9812 12336
rect 9673 12278 9812 12280
rect 9673 12275 9739 12278
rect 9806 12276 9812 12278
rect 9876 12276 9882 12340
rect 9952 12338 10012 12550
rect 10816 12544 11132 12545
rect 10816 12480 10822 12544
rect 10886 12480 10902 12544
rect 10966 12480 10982 12544
rect 11046 12480 11062 12544
rect 11126 12480 11132 12544
rect 10816 12479 11132 12480
rect 14764 12544 15080 12545
rect 14764 12480 14770 12544
rect 14834 12480 14850 12544
rect 14914 12480 14930 12544
rect 14994 12480 15010 12544
rect 15074 12480 15080 12544
rect 14764 12479 15080 12480
rect 10777 12338 10843 12341
rect 9952 12336 10843 12338
rect 9952 12280 10782 12336
rect 10838 12280 10843 12336
rect 9952 12278 10843 12280
rect 10777 12275 10843 12278
rect 6821 12202 6887 12205
rect 11513 12202 11579 12205
rect 6821 12200 11579 12202
rect 6821 12144 6826 12200
rect 6882 12144 11518 12200
rect 11574 12144 11579 12200
rect 6821 12142 11579 12144
rect 6821 12139 6887 12142
rect 11513 12139 11579 12142
rect 8569 12068 8635 12069
rect 8518 12004 8524 12068
rect 8588 12066 8635 12068
rect 8588 12064 8680 12066
rect 8630 12008 8680 12064
rect 8588 12006 8680 12008
rect 8588 12004 8635 12006
rect 9254 12004 9260 12068
rect 9324 12066 9330 12068
rect 9581 12066 9647 12069
rect 9324 12064 9647 12066
rect 9324 12008 9586 12064
rect 9642 12008 9647 12064
rect 9324 12006 9647 12008
rect 9324 12004 9330 12006
rect 8569 12003 8635 12004
rect 9581 12003 9647 12006
rect 4894 12000 5210 12001
rect 4894 11936 4900 12000
rect 4964 11936 4980 12000
rect 5044 11936 5060 12000
rect 5124 11936 5140 12000
rect 5204 11936 5210 12000
rect 4894 11935 5210 11936
rect 8842 12000 9158 12001
rect 8842 11936 8848 12000
rect 8912 11936 8928 12000
rect 8992 11936 9008 12000
rect 9072 11936 9088 12000
rect 9152 11936 9158 12000
rect 8842 11935 9158 11936
rect 12790 12000 13106 12001
rect 12790 11936 12796 12000
rect 12860 11936 12876 12000
rect 12940 11936 12956 12000
rect 13020 11936 13036 12000
rect 13100 11936 13106 12000
rect 12790 11935 13106 11936
rect 3550 11732 3556 11796
rect 3620 11794 3626 11796
rect 7925 11794 7991 11797
rect 8201 11794 8267 11797
rect 3620 11792 8267 11794
rect 3620 11736 7930 11792
rect 7986 11736 8206 11792
rect 8262 11736 8267 11792
rect 3620 11734 8267 11736
rect 3620 11732 3626 11734
rect 7925 11731 7991 11734
rect 8201 11731 8267 11734
rect 8702 11732 8708 11796
rect 8772 11794 8778 11796
rect 9397 11794 9463 11797
rect 8772 11792 9463 11794
rect 8772 11736 9402 11792
rect 9458 11736 9463 11792
rect 8772 11734 9463 11736
rect 8772 11732 8778 11734
rect 9397 11731 9463 11734
rect 10542 11732 10548 11796
rect 10612 11794 10618 11796
rect 10685 11794 10751 11797
rect 13905 11794 13971 11797
rect 10612 11792 13971 11794
rect 10612 11736 10690 11792
rect 10746 11736 13910 11792
rect 13966 11736 13971 11792
rect 10612 11734 13971 11736
rect 10612 11732 10618 11734
rect 10685 11731 10751 11734
rect 13905 11731 13971 11734
rect 4245 11658 4311 11661
rect 7465 11658 7531 11661
rect 7833 11658 7899 11661
rect 10133 11658 10199 11661
rect 4245 11656 7712 11658
rect 4245 11600 4250 11656
rect 4306 11600 7470 11656
rect 7526 11600 7712 11656
rect 4245 11598 7712 11600
rect 4245 11595 4311 11598
rect 7465 11595 7531 11598
rect 3734 11460 3740 11524
rect 3804 11522 3810 11524
rect 6637 11522 6703 11525
rect 3804 11520 6703 11522
rect 3804 11464 6642 11520
rect 6698 11464 6703 11520
rect 3804 11462 6703 11464
rect 7652 11522 7712 11598
rect 7833 11656 10199 11658
rect 7833 11600 7838 11656
rect 7894 11600 10138 11656
rect 10194 11600 10199 11656
rect 7833 11598 10199 11600
rect 7833 11595 7899 11598
rect 10133 11595 10199 11598
rect 9121 11522 9187 11525
rect 7652 11520 9187 11522
rect 7652 11464 9126 11520
rect 9182 11464 9187 11520
rect 7652 11462 9187 11464
rect 3804 11460 3810 11462
rect 6637 11459 6703 11462
rect 9121 11459 9187 11462
rect 9673 11522 9739 11525
rect 10501 11522 10567 11525
rect 9673 11520 10567 11522
rect 9673 11464 9678 11520
rect 9734 11464 10506 11520
rect 10562 11464 10567 11520
rect 9673 11462 10567 11464
rect 9673 11459 9739 11462
rect 10501 11459 10567 11462
rect 2920 11456 3236 11457
rect 2920 11392 2926 11456
rect 2990 11392 3006 11456
rect 3070 11392 3086 11456
rect 3150 11392 3166 11456
rect 3230 11392 3236 11456
rect 2920 11391 3236 11392
rect 6868 11456 7184 11457
rect 6868 11392 6874 11456
rect 6938 11392 6954 11456
rect 7018 11392 7034 11456
rect 7098 11392 7114 11456
rect 7178 11392 7184 11456
rect 6868 11391 7184 11392
rect 10816 11456 11132 11457
rect 10816 11392 10822 11456
rect 10886 11392 10902 11456
rect 10966 11392 10982 11456
rect 11046 11392 11062 11456
rect 11126 11392 11132 11456
rect 10816 11391 11132 11392
rect 14764 11456 15080 11457
rect 14764 11392 14770 11456
rect 14834 11392 14850 11456
rect 14914 11392 14930 11456
rect 14994 11392 15010 11456
rect 15074 11392 15080 11456
rect 14764 11391 15080 11392
rect 0 11160 400 11280
rect 7833 11250 7899 11253
rect 5766 11248 7899 11250
rect 5766 11192 7838 11248
rect 7894 11192 7899 11248
rect 5766 11190 7899 11192
rect 2630 11052 2636 11116
rect 2700 11114 2706 11116
rect 5766 11114 5826 11190
rect 7833 11187 7899 11190
rect 8845 11250 8911 11253
rect 10133 11250 10199 11253
rect 8845 11248 10199 11250
rect 8845 11192 8850 11248
rect 8906 11192 10138 11248
rect 10194 11192 10199 11248
rect 8845 11190 10199 11192
rect 8845 11187 8911 11190
rect 10133 11187 10199 11190
rect 11145 11250 11211 11253
rect 12433 11250 12499 11253
rect 11145 11248 12499 11250
rect 11145 11192 11150 11248
rect 11206 11192 12438 11248
rect 12494 11192 12499 11248
rect 11145 11190 12499 11192
rect 11145 11187 11211 11190
rect 12433 11187 12499 11190
rect 2700 11054 5826 11114
rect 2700 11052 2706 11054
rect 5942 11052 5948 11116
rect 6012 11114 6018 11116
rect 9029 11114 9095 11117
rect 6012 11112 9095 11114
rect 6012 11056 9034 11112
rect 9090 11056 9095 11112
rect 6012 11054 9095 11056
rect 6012 11052 6018 11054
rect 9029 11051 9095 11054
rect 9213 11114 9279 11117
rect 10777 11114 10843 11117
rect 13445 11114 13511 11117
rect 9213 11112 9920 11114
rect 9213 11056 9218 11112
rect 9274 11056 9920 11112
rect 9213 11054 9920 11056
rect 9213 11051 9279 11054
rect 9860 10978 9920 11054
rect 10777 11112 13511 11114
rect 10777 11056 10782 11112
rect 10838 11056 13450 11112
rect 13506 11056 13511 11112
rect 10777 11054 13511 11056
rect 10777 11051 10843 11054
rect 13445 11051 13511 11054
rect 12065 10978 12131 10981
rect 9860 10976 12131 10978
rect 9860 10920 12070 10976
rect 12126 10920 12131 10976
rect 9860 10918 12131 10920
rect 12065 10915 12131 10918
rect 4894 10912 5210 10913
rect 4894 10848 4900 10912
rect 4964 10848 4980 10912
rect 5044 10848 5060 10912
rect 5124 10848 5140 10912
rect 5204 10848 5210 10912
rect 4894 10847 5210 10848
rect 8842 10912 9158 10913
rect 8842 10848 8848 10912
rect 8912 10848 8928 10912
rect 8992 10848 9008 10912
rect 9072 10848 9088 10912
rect 9152 10848 9158 10912
rect 8842 10847 9158 10848
rect 12790 10912 13106 10913
rect 12790 10848 12796 10912
rect 12860 10848 12876 10912
rect 12940 10848 12956 10912
rect 13020 10848 13036 10912
rect 13100 10848 13106 10912
rect 12790 10847 13106 10848
rect 9673 10842 9739 10845
rect 9806 10842 9812 10844
rect 9673 10840 9812 10842
rect 9673 10784 9678 10840
rect 9734 10784 9812 10840
rect 9673 10782 9812 10784
rect 9673 10779 9739 10782
rect 9806 10780 9812 10782
rect 9876 10842 9882 10844
rect 10869 10842 10935 10845
rect 11697 10842 11763 10845
rect 9876 10840 11763 10842
rect 9876 10784 10874 10840
rect 10930 10784 11702 10840
rect 11758 10784 11763 10840
rect 9876 10782 11763 10784
rect 9876 10780 9882 10782
rect 10869 10779 10935 10782
rect 11697 10779 11763 10782
rect 2773 10706 2839 10709
rect 5625 10706 5691 10709
rect 2773 10704 5691 10706
rect 2773 10648 2778 10704
rect 2834 10648 5630 10704
rect 5686 10648 5691 10704
rect 2773 10646 5691 10648
rect 2773 10643 2839 10646
rect 5625 10643 5691 10646
rect 8150 10644 8156 10708
rect 8220 10706 8226 10708
rect 8753 10706 8819 10709
rect 8220 10704 8819 10706
rect 8220 10648 8758 10704
rect 8814 10648 8819 10704
rect 8220 10646 8819 10648
rect 8220 10644 8226 10646
rect 8753 10643 8819 10646
rect 8937 10706 9003 10709
rect 13813 10706 13879 10709
rect 8937 10704 13879 10706
rect 8937 10648 8942 10704
rect 8998 10648 13818 10704
rect 13874 10648 13879 10704
rect 8937 10646 13879 10648
rect 8937 10643 9003 10646
rect 13813 10643 13879 10646
rect 2497 10570 2563 10573
rect 11145 10570 11211 10573
rect 2497 10568 11211 10570
rect 2497 10512 2502 10568
rect 2558 10512 11150 10568
rect 11206 10512 11211 10568
rect 2497 10510 11211 10512
rect 2497 10507 2563 10510
rect 11145 10507 11211 10510
rect 7966 10372 7972 10436
rect 8036 10434 8042 10436
rect 9857 10434 9923 10437
rect 8036 10432 10426 10434
rect 8036 10376 9862 10432
rect 9918 10376 10426 10432
rect 8036 10374 10426 10376
rect 8036 10372 8042 10374
rect 9857 10371 9923 10374
rect 2920 10368 3236 10369
rect 2920 10304 2926 10368
rect 2990 10304 3006 10368
rect 3070 10304 3086 10368
rect 3150 10304 3166 10368
rect 3230 10304 3236 10368
rect 2920 10303 3236 10304
rect 6868 10368 7184 10369
rect 6868 10304 6874 10368
rect 6938 10304 6954 10368
rect 7018 10304 7034 10368
rect 7098 10304 7114 10368
rect 7178 10304 7184 10368
rect 6868 10303 7184 10304
rect 7414 10236 7420 10300
rect 7484 10298 7490 10300
rect 7649 10298 7715 10301
rect 8937 10298 9003 10301
rect 7484 10296 9003 10298
rect 7484 10240 7654 10296
rect 7710 10240 8942 10296
rect 8998 10240 9003 10296
rect 7484 10238 9003 10240
rect 10366 10298 10426 10374
rect 10816 10368 11132 10369
rect 10816 10304 10822 10368
rect 10886 10304 10902 10368
rect 10966 10304 10982 10368
rect 11046 10304 11062 10368
rect 11126 10304 11132 10368
rect 10816 10303 11132 10304
rect 14764 10368 15080 10369
rect 14764 10304 14770 10368
rect 14834 10304 14850 10368
rect 14914 10304 14930 10368
rect 14994 10304 15010 10368
rect 15074 10304 15080 10368
rect 14764 10303 15080 10304
rect 10685 10298 10751 10301
rect 10366 10296 10751 10298
rect 10366 10240 10690 10296
rect 10746 10240 10751 10296
rect 10366 10238 10751 10240
rect 7484 10236 7490 10238
rect 7649 10235 7715 10238
rect 8937 10235 9003 10238
rect 10685 10235 10751 10238
rect 3417 10162 3483 10165
rect 14457 10162 14523 10165
rect 3417 10160 14523 10162
rect 3417 10104 3422 10160
rect 3478 10104 14462 10160
rect 14518 10104 14523 10160
rect 3417 10102 14523 10104
rect 3417 10099 3483 10102
rect 14457 10099 14523 10102
rect 1761 10026 1827 10029
rect 2630 10026 2636 10028
rect 1761 10024 2636 10026
rect 1761 9968 1766 10024
rect 1822 9968 2636 10024
rect 1761 9966 2636 9968
rect 1761 9963 1827 9966
rect 2630 9964 2636 9966
rect 2700 9964 2706 10028
rect 4061 10026 4127 10029
rect 11881 10026 11947 10029
rect 4061 10024 11947 10026
rect 4061 9968 4066 10024
rect 4122 9968 11886 10024
rect 11942 9968 11947 10024
rect 4061 9966 11947 9968
rect 4061 9963 4127 9966
rect 11881 9963 11947 9966
rect 9581 9890 9647 9893
rect 11789 9890 11855 9893
rect 9581 9888 11855 9890
rect 9581 9832 9586 9888
rect 9642 9832 11794 9888
rect 11850 9832 11855 9888
rect 9581 9830 11855 9832
rect 9581 9827 9647 9830
rect 11789 9827 11855 9830
rect 4894 9824 5210 9825
rect 0 9664 400 9784
rect 4894 9760 4900 9824
rect 4964 9760 4980 9824
rect 5044 9760 5060 9824
rect 5124 9760 5140 9824
rect 5204 9760 5210 9824
rect 4894 9759 5210 9760
rect 8842 9824 9158 9825
rect 8842 9760 8848 9824
rect 8912 9760 8928 9824
rect 8992 9760 9008 9824
rect 9072 9760 9088 9824
rect 9152 9760 9158 9824
rect 8842 9759 9158 9760
rect 12790 9824 13106 9825
rect 12790 9760 12796 9824
rect 12860 9760 12876 9824
rect 12940 9760 12956 9824
rect 13020 9760 13036 9824
rect 13100 9760 13106 9824
rect 12790 9759 13106 9760
rect 9622 9692 9628 9756
rect 9692 9754 9698 9756
rect 10041 9754 10107 9757
rect 9692 9752 10107 9754
rect 9692 9696 10046 9752
rect 10102 9696 10107 9752
rect 9692 9694 10107 9696
rect 9692 9692 9698 9694
rect 10041 9691 10107 9694
rect 4654 9556 4660 9620
rect 4724 9618 4730 9620
rect 12341 9618 12407 9621
rect 4724 9616 12407 9618
rect 4724 9560 12346 9616
rect 12402 9560 12407 9616
rect 4724 9558 12407 9560
rect 4724 9556 4730 9558
rect 12341 9555 12407 9558
rect 1301 9482 1367 9485
rect 8201 9482 8267 9485
rect 9949 9484 10015 9485
rect 9949 9482 9996 9484
rect 1301 9480 8267 9482
rect 1301 9424 1306 9480
rect 1362 9424 8206 9480
rect 8262 9424 8267 9480
rect 1301 9422 8267 9424
rect 9904 9480 9996 9482
rect 9904 9424 9954 9480
rect 9904 9422 9996 9424
rect 1301 9419 1367 9422
rect 8201 9419 8267 9422
rect 9949 9420 9996 9422
rect 10060 9420 10066 9484
rect 12433 9482 12499 9485
rect 10688 9480 12499 9482
rect 10688 9424 12438 9480
rect 12494 9424 12499 9480
rect 10688 9422 12499 9424
rect 9949 9419 10015 9420
rect 7649 9346 7715 9349
rect 8201 9346 8267 9349
rect 7649 9344 8267 9346
rect 7649 9288 7654 9344
rect 7710 9288 8206 9344
rect 8262 9288 8267 9344
rect 7649 9286 8267 9288
rect 7649 9283 7715 9286
rect 8201 9283 8267 9286
rect 8569 9346 8635 9349
rect 9397 9346 9463 9349
rect 8569 9344 9463 9346
rect 8569 9288 8574 9344
rect 8630 9288 9402 9344
rect 9458 9288 9463 9344
rect 8569 9286 9463 9288
rect 8569 9283 8635 9286
rect 9397 9283 9463 9286
rect 10133 9346 10199 9349
rect 10688 9346 10748 9422
rect 12433 9419 12499 9422
rect 10133 9344 10748 9346
rect 10133 9288 10138 9344
rect 10194 9288 10748 9344
rect 10133 9286 10748 9288
rect 10133 9283 10199 9286
rect 2920 9280 3236 9281
rect 2920 9216 2926 9280
rect 2990 9216 3006 9280
rect 3070 9216 3086 9280
rect 3150 9216 3166 9280
rect 3230 9216 3236 9280
rect 2920 9215 3236 9216
rect 6868 9280 7184 9281
rect 6868 9216 6874 9280
rect 6938 9216 6954 9280
rect 7018 9216 7034 9280
rect 7098 9216 7114 9280
rect 7178 9216 7184 9280
rect 6868 9215 7184 9216
rect 10816 9280 11132 9281
rect 10816 9216 10822 9280
rect 10886 9216 10902 9280
rect 10966 9216 10982 9280
rect 11046 9216 11062 9280
rect 11126 9216 11132 9280
rect 10816 9215 11132 9216
rect 14764 9280 15080 9281
rect 14764 9216 14770 9280
rect 14834 9216 14850 9280
rect 14914 9216 14930 9280
rect 14994 9216 15010 9280
rect 15074 9216 15080 9280
rect 14764 9215 15080 9216
rect 7649 9210 7715 9213
rect 9254 9210 9260 9212
rect 7649 9208 9260 9210
rect 7649 9152 7654 9208
rect 7710 9152 9260 9208
rect 7649 9150 9260 9152
rect 7649 9147 7715 9150
rect 9254 9148 9260 9150
rect 9324 9148 9330 9212
rect 9673 9210 9739 9213
rect 10174 9210 10180 9212
rect 9673 9208 10180 9210
rect 9673 9152 9678 9208
rect 9734 9152 10180 9208
rect 9673 9150 10180 9152
rect 9673 9147 9739 9150
rect 10174 9148 10180 9150
rect 10244 9148 10250 9212
rect 10358 9148 10364 9212
rect 10428 9210 10434 9212
rect 10501 9210 10567 9213
rect 10428 9208 10567 9210
rect 10428 9152 10506 9208
rect 10562 9152 10567 9208
rect 10428 9150 10567 9152
rect 10428 9148 10434 9150
rect 10501 9147 10567 9150
rect 1485 9074 1551 9077
rect 6545 9074 6611 9077
rect 8017 9074 8083 9077
rect 1485 9072 8083 9074
rect 1485 9016 1490 9072
rect 1546 9016 6550 9072
rect 6606 9016 8022 9072
rect 8078 9016 8083 9072
rect 1485 9014 8083 9016
rect 1485 9011 1551 9014
rect 6545 9011 6611 9014
rect 8017 9011 8083 9014
rect 8661 9074 8727 9077
rect 9857 9074 9923 9077
rect 8661 9072 9923 9074
rect 8661 9016 8666 9072
rect 8722 9016 9862 9072
rect 9918 9016 9923 9072
rect 8661 9014 9923 9016
rect 8661 9011 8727 9014
rect 9857 9011 9923 9014
rect 11789 9074 11855 9077
rect 11973 9074 12039 9077
rect 11789 9072 12039 9074
rect 11789 9016 11794 9072
rect 11850 9016 11978 9072
rect 12034 9016 12039 9072
rect 11789 9014 12039 9016
rect 11789 9011 11855 9014
rect 11973 9011 12039 9014
rect 3509 8938 3575 8941
rect 6085 8938 6151 8941
rect 3509 8936 6151 8938
rect 3509 8880 3514 8936
rect 3570 8880 6090 8936
rect 6146 8880 6151 8936
rect 3509 8878 6151 8880
rect 3509 8875 3575 8878
rect 6085 8875 6151 8878
rect 7097 8938 7163 8941
rect 8334 8938 8340 8940
rect 7097 8936 8340 8938
rect 7097 8880 7102 8936
rect 7158 8880 8340 8936
rect 7097 8878 8340 8880
rect 7097 8875 7163 8878
rect 8334 8876 8340 8878
rect 8404 8938 8410 8940
rect 11053 8938 11119 8941
rect 8404 8936 11119 8938
rect 8404 8880 11058 8936
rect 11114 8880 11119 8936
rect 8404 8878 11119 8880
rect 8404 8876 8410 8878
rect 11053 8875 11119 8878
rect 11237 8936 11303 8941
rect 11237 8880 11242 8936
rect 11298 8880 11303 8936
rect 11237 8875 11303 8880
rect 6678 8740 6684 8804
rect 6748 8802 6754 8804
rect 8201 8802 8267 8805
rect 6748 8800 8267 8802
rect 6748 8744 8206 8800
rect 8262 8744 8267 8800
rect 6748 8742 8267 8744
rect 6748 8740 6754 8742
rect 8201 8739 8267 8742
rect 9438 8740 9444 8804
rect 9508 8802 9514 8804
rect 10593 8802 10659 8805
rect 9508 8800 10659 8802
rect 9508 8744 10598 8800
rect 10654 8744 10659 8800
rect 9508 8742 10659 8744
rect 9508 8740 9514 8742
rect 10593 8739 10659 8742
rect 10777 8802 10843 8805
rect 11240 8802 11300 8875
rect 10777 8800 11300 8802
rect 10777 8744 10782 8800
rect 10838 8744 11300 8800
rect 10777 8742 11300 8744
rect 10777 8739 10843 8742
rect 4894 8736 5210 8737
rect 4894 8672 4900 8736
rect 4964 8672 4980 8736
rect 5044 8672 5060 8736
rect 5124 8672 5140 8736
rect 5204 8672 5210 8736
rect 4894 8671 5210 8672
rect 8842 8736 9158 8737
rect 8842 8672 8848 8736
rect 8912 8672 8928 8736
rect 8992 8672 9008 8736
rect 9072 8672 9088 8736
rect 9152 8672 9158 8736
rect 8842 8671 9158 8672
rect 12790 8736 13106 8737
rect 12790 8672 12796 8736
rect 12860 8672 12876 8736
rect 12940 8672 12956 8736
rect 13020 8672 13036 8736
rect 13100 8672 13106 8736
rect 12790 8671 13106 8672
rect 8569 8666 8635 8669
rect 5398 8664 8635 8666
rect 5398 8608 8574 8664
rect 8630 8608 8635 8664
rect 5398 8606 8635 8608
rect 2681 8530 2747 8533
rect 4705 8530 4771 8533
rect 2681 8528 4771 8530
rect 2681 8472 2686 8528
rect 2742 8472 4710 8528
rect 4766 8472 4771 8528
rect 2681 8470 4771 8472
rect 2681 8467 2747 8470
rect 4705 8467 4771 8470
rect 5073 8530 5139 8533
rect 5398 8530 5458 8606
rect 8569 8603 8635 8606
rect 9254 8604 9260 8668
rect 9324 8666 9330 8668
rect 10869 8666 10935 8669
rect 9324 8664 10935 8666
rect 9324 8608 10874 8664
rect 10930 8608 10935 8664
rect 9324 8606 10935 8608
rect 9324 8604 9330 8606
rect 10869 8603 10935 8606
rect 5073 8528 5458 8530
rect 5073 8472 5078 8528
rect 5134 8472 5458 8528
rect 5073 8470 5458 8472
rect 6821 8530 6887 8533
rect 12157 8530 12223 8533
rect 6821 8528 12223 8530
rect 6821 8472 6826 8528
rect 6882 8472 12162 8528
rect 12218 8472 12223 8528
rect 6821 8470 12223 8472
rect 5073 8467 5139 8470
rect 6821 8467 6887 8470
rect 12157 8467 12223 8470
rect 3509 8394 3575 8397
rect 5574 8394 5580 8396
rect 3509 8392 5580 8394
rect 3509 8336 3514 8392
rect 3570 8336 5580 8392
rect 3509 8334 5580 8336
rect 3509 8331 3575 8334
rect 5574 8332 5580 8334
rect 5644 8332 5650 8396
rect 6686 8334 7344 8394
rect 0 8258 400 8288
rect 3969 8258 4035 8261
rect 6686 8258 6746 8334
rect 0 8198 2790 8258
rect 0 8168 400 8198
rect 2730 7986 2790 8198
rect 3969 8256 6746 8258
rect 3969 8200 3974 8256
rect 4030 8200 6746 8256
rect 3969 8198 6746 8200
rect 7284 8258 7344 8334
rect 7414 8332 7420 8396
rect 7484 8394 7490 8396
rect 7557 8394 7623 8397
rect 7484 8392 7623 8394
rect 7484 8336 7562 8392
rect 7618 8336 7623 8392
rect 7484 8334 7623 8336
rect 7484 8332 7490 8334
rect 7557 8331 7623 8334
rect 8702 8332 8708 8396
rect 8772 8394 8778 8396
rect 9029 8394 9095 8397
rect 9438 8394 9444 8396
rect 8772 8392 9444 8394
rect 8772 8336 9034 8392
rect 9090 8336 9444 8392
rect 8772 8334 9444 8336
rect 8772 8332 8778 8334
rect 9029 8331 9095 8334
rect 9438 8332 9444 8334
rect 9508 8332 9514 8396
rect 9806 8332 9812 8396
rect 9876 8394 9882 8396
rect 10041 8394 10107 8397
rect 9876 8392 10107 8394
rect 9876 8336 10046 8392
rect 10102 8336 10107 8392
rect 9876 8334 10107 8336
rect 9876 8332 9882 8334
rect 10041 8331 10107 8334
rect 11237 8396 11303 8397
rect 11237 8392 11284 8396
rect 11348 8394 11354 8396
rect 11237 8336 11242 8392
rect 11237 8332 11284 8336
rect 11348 8334 11394 8394
rect 11348 8332 11354 8334
rect 11237 8331 11303 8332
rect 10409 8258 10475 8261
rect 7284 8256 10475 8258
rect 7284 8200 10414 8256
rect 10470 8200 10475 8256
rect 7284 8198 10475 8200
rect 3969 8195 4035 8198
rect 10409 8195 10475 8198
rect 2920 8192 3236 8193
rect 2920 8128 2926 8192
rect 2990 8128 3006 8192
rect 3070 8128 3086 8192
rect 3150 8128 3166 8192
rect 3230 8128 3236 8192
rect 2920 8127 3236 8128
rect 6868 8192 7184 8193
rect 6868 8128 6874 8192
rect 6938 8128 6954 8192
rect 7018 8128 7034 8192
rect 7098 8128 7114 8192
rect 7178 8128 7184 8192
rect 6868 8127 7184 8128
rect 10816 8192 11132 8193
rect 10816 8128 10822 8192
rect 10886 8128 10902 8192
rect 10966 8128 10982 8192
rect 11046 8128 11062 8192
rect 11126 8128 11132 8192
rect 10816 8127 11132 8128
rect 14764 8192 15080 8193
rect 14764 8128 14770 8192
rect 14834 8128 14850 8192
rect 14914 8128 14930 8192
rect 14994 8128 15010 8192
rect 15074 8128 15080 8192
rect 14764 8127 15080 8128
rect 5717 8124 5783 8125
rect 6177 8124 6243 8125
rect 6361 8124 6427 8125
rect 5717 8120 5764 8124
rect 5828 8122 5834 8124
rect 6126 8122 6132 8124
rect 5717 8064 5722 8120
rect 5717 8060 5764 8064
rect 5828 8062 5874 8122
rect 6086 8062 6132 8122
rect 6196 8120 6243 8124
rect 6238 8064 6243 8120
rect 5828 8060 5834 8062
rect 6126 8060 6132 8062
rect 6196 8060 6243 8064
rect 6310 8060 6316 8124
rect 6380 8122 6427 8124
rect 8937 8122 9003 8125
rect 10542 8122 10548 8124
rect 6380 8120 6472 8122
rect 6422 8064 6472 8120
rect 6380 8062 6472 8064
rect 8937 8120 10548 8122
rect 8937 8064 8942 8120
rect 8998 8064 10548 8120
rect 8937 8062 10548 8064
rect 6380 8060 6427 8062
rect 5717 8059 5783 8060
rect 6177 8059 6243 8060
rect 6361 8059 6427 8060
rect 8937 8059 9003 8062
rect 10542 8060 10548 8062
rect 10612 8060 10618 8124
rect 3417 7986 3483 7989
rect 2730 7984 3483 7986
rect 2730 7928 3422 7984
rect 3478 7928 3483 7984
rect 2730 7926 3483 7928
rect 3417 7923 3483 7926
rect 4705 7986 4771 7989
rect 6361 7986 6427 7989
rect 4705 7984 6427 7986
rect 4705 7928 4710 7984
rect 4766 7928 6366 7984
rect 6422 7928 6427 7984
rect 4705 7926 6427 7928
rect 4705 7923 4771 7926
rect 6361 7923 6427 7926
rect 7097 7986 7163 7989
rect 13537 7986 13603 7989
rect 7097 7984 13603 7986
rect 7097 7928 7102 7984
rect 7158 7928 13542 7984
rect 13598 7928 13603 7984
rect 7097 7926 13603 7928
rect 7097 7923 7163 7926
rect 13537 7923 13603 7926
rect 2037 7850 2103 7853
rect 7465 7850 7531 7853
rect 10358 7850 10364 7852
rect 2037 7848 7531 7850
rect 2037 7792 2042 7848
rect 2098 7792 7470 7848
rect 7526 7792 7531 7848
rect 2037 7790 7531 7792
rect 2037 7787 2103 7790
rect 7465 7787 7531 7790
rect 8388 7790 10364 7850
rect 8388 7717 8448 7790
rect 10358 7788 10364 7790
rect 10428 7788 10434 7852
rect 5533 7714 5599 7717
rect 5533 7712 7896 7714
rect 5533 7656 5538 7712
rect 5594 7656 7896 7712
rect 5533 7654 7896 7656
rect 5533 7651 5599 7654
rect 4894 7648 5210 7649
rect 4894 7584 4900 7648
rect 4964 7584 4980 7648
rect 5044 7584 5060 7648
rect 5124 7584 5140 7648
rect 5204 7584 5210 7648
rect 4894 7583 5210 7584
rect 7836 7581 7896 7654
rect 8385 7712 8451 7717
rect 8385 7656 8390 7712
rect 8446 7656 8451 7712
rect 8385 7651 8451 7656
rect 9673 7714 9739 7717
rect 10174 7714 10180 7716
rect 9673 7712 10180 7714
rect 9673 7656 9678 7712
rect 9734 7656 10180 7712
rect 9673 7654 10180 7656
rect 9673 7651 9739 7654
rect 10174 7652 10180 7654
rect 10244 7652 10250 7716
rect 8842 7648 9158 7649
rect 8842 7584 8848 7648
rect 8912 7584 8928 7648
rect 8992 7584 9008 7648
rect 9072 7584 9088 7648
rect 9152 7584 9158 7648
rect 8842 7583 9158 7584
rect 12790 7648 13106 7649
rect 12790 7584 12796 7648
rect 12860 7584 12876 7648
rect 12940 7584 12956 7648
rect 13020 7584 13036 7648
rect 13100 7584 13106 7648
rect 12790 7583 13106 7584
rect 5901 7580 5967 7581
rect 5901 7576 5948 7580
rect 6012 7578 6018 7580
rect 7097 7578 7163 7581
rect 5901 7520 5906 7576
rect 5901 7516 5948 7520
rect 6012 7518 6058 7578
rect 6686 7576 7163 7578
rect 6686 7520 7102 7576
rect 7158 7520 7163 7576
rect 6686 7518 7163 7520
rect 6012 7516 6018 7518
rect 5901 7515 5967 7516
rect 4245 7442 4311 7445
rect 6686 7442 6746 7518
rect 7097 7515 7163 7518
rect 7833 7576 7899 7581
rect 7833 7520 7838 7576
rect 7894 7520 7899 7576
rect 7833 7515 7899 7520
rect 9857 7578 9923 7581
rect 9990 7578 9996 7580
rect 9857 7576 9996 7578
rect 9857 7520 9862 7576
rect 9918 7520 9996 7576
rect 9857 7518 9996 7520
rect 9857 7515 9923 7518
rect 9990 7516 9996 7518
rect 10060 7516 10066 7580
rect 4245 7440 6746 7442
rect 4245 7384 4250 7440
rect 4306 7384 6746 7440
rect 4245 7382 6746 7384
rect 6821 7442 6887 7445
rect 9029 7442 9095 7445
rect 6821 7440 9095 7442
rect 6821 7384 6826 7440
rect 6882 7384 9034 7440
rect 9090 7384 9095 7440
rect 6821 7382 9095 7384
rect 4245 7379 4311 7382
rect 6821 7379 6887 7382
rect 9029 7379 9095 7382
rect 1853 7306 1919 7309
rect 9397 7306 9463 7309
rect 12525 7306 12591 7309
rect 1853 7304 9463 7306
rect 1853 7248 1858 7304
rect 1914 7248 9402 7304
rect 9458 7248 9463 7304
rect 1853 7246 9463 7248
rect 1853 7243 1919 7246
rect 9397 7243 9463 7246
rect 9630 7304 12591 7306
rect 9630 7248 12530 7304
rect 12586 7248 12591 7304
rect 9630 7246 12591 7248
rect 5625 7170 5691 7173
rect 6126 7170 6132 7172
rect 5625 7168 6132 7170
rect 5625 7112 5630 7168
rect 5686 7112 6132 7168
rect 5625 7110 6132 7112
rect 5625 7107 5691 7110
rect 6126 7108 6132 7110
rect 6196 7108 6202 7172
rect 6361 7170 6427 7173
rect 6494 7170 6500 7172
rect 6361 7168 6500 7170
rect 6361 7112 6366 7168
rect 6422 7112 6500 7168
rect 6361 7110 6500 7112
rect 6361 7107 6427 7110
rect 6494 7108 6500 7110
rect 6564 7108 6570 7172
rect 7833 7170 7899 7173
rect 9397 7170 9463 7173
rect 7833 7168 9463 7170
rect 7833 7112 7838 7168
rect 7894 7112 9402 7168
rect 9458 7112 9463 7168
rect 7833 7110 9463 7112
rect 7833 7107 7899 7110
rect 9397 7107 9463 7110
rect 2920 7104 3236 7105
rect 2920 7040 2926 7104
rect 2990 7040 3006 7104
rect 3070 7040 3086 7104
rect 3150 7040 3166 7104
rect 3230 7040 3236 7104
rect 2920 7039 3236 7040
rect 6868 7104 7184 7105
rect 6868 7040 6874 7104
rect 6938 7040 6954 7104
rect 7018 7040 7034 7104
rect 7098 7040 7114 7104
rect 7178 7040 7184 7104
rect 6868 7039 7184 7040
rect 4153 7036 4219 7037
rect 4102 7034 4108 7036
rect 4062 6974 4108 7034
rect 4172 7032 4219 7036
rect 4214 6976 4219 7032
rect 4102 6972 4108 6974
rect 4172 6972 4219 6976
rect 4153 6971 4219 6972
rect 5165 7034 5231 7037
rect 9630 7034 9690 7246
rect 12525 7243 12591 7246
rect 10816 7104 11132 7105
rect 10816 7040 10822 7104
rect 10886 7040 10902 7104
rect 10966 7040 10982 7104
rect 11046 7040 11062 7104
rect 11126 7040 11132 7104
rect 10816 7039 11132 7040
rect 14764 7104 15080 7105
rect 14764 7040 14770 7104
rect 14834 7040 14850 7104
rect 14914 7040 14930 7104
rect 14994 7040 15010 7104
rect 15074 7040 15080 7104
rect 14764 7039 15080 7040
rect 5165 7032 6746 7034
rect 5165 6976 5170 7032
rect 5226 6976 6746 7032
rect 5165 6974 6746 6976
rect 5165 6971 5231 6974
rect 4061 6898 4127 6901
rect 5625 6898 5691 6901
rect 6361 6900 6427 6901
rect 4061 6896 5691 6898
rect 4061 6840 4066 6896
rect 4122 6840 5630 6896
rect 5686 6840 5691 6896
rect 4061 6838 5691 6840
rect 4061 6835 4127 6838
rect 5625 6835 5691 6838
rect 6310 6836 6316 6900
rect 6380 6898 6427 6900
rect 6686 6898 6746 6974
rect 7284 6974 9690 7034
rect 7284 6901 7344 6974
rect 7281 6898 7347 6901
rect 6380 6896 6472 6898
rect 6422 6840 6472 6896
rect 6380 6838 6472 6840
rect 6686 6896 7347 6898
rect 6686 6840 7286 6896
rect 7342 6840 7347 6896
rect 6686 6838 7347 6840
rect 6380 6836 6427 6838
rect 6361 6835 6427 6836
rect 7281 6835 7347 6838
rect 7557 6898 7623 6901
rect 10317 6898 10383 6901
rect 7557 6896 10383 6898
rect 7557 6840 7562 6896
rect 7618 6840 10322 6896
rect 10378 6840 10383 6896
rect 7557 6838 10383 6840
rect 7557 6835 7623 6838
rect 10317 6835 10383 6838
rect 0 6762 400 6792
rect 1393 6762 1459 6765
rect 0 6760 1459 6762
rect 0 6704 1398 6760
rect 1454 6704 1459 6760
rect 0 6702 1459 6704
rect 0 6672 400 6702
rect 1393 6699 1459 6702
rect 4705 6762 4771 6765
rect 12709 6762 12775 6765
rect 4705 6760 12775 6762
rect 4705 6704 4710 6760
rect 4766 6704 12714 6760
rect 12770 6704 12775 6760
rect 4705 6702 12775 6704
rect 4705 6699 4771 6702
rect 12709 6699 12775 6702
rect 5809 6628 5875 6629
rect 5758 6564 5764 6628
rect 5828 6626 5875 6628
rect 6085 6626 6151 6629
rect 8150 6626 8156 6628
rect 5828 6624 5920 6626
rect 5870 6568 5920 6624
rect 5828 6566 5920 6568
rect 6085 6624 8156 6626
rect 6085 6568 6090 6624
rect 6146 6568 8156 6624
rect 6085 6566 8156 6568
rect 5828 6564 5875 6566
rect 5809 6563 5875 6564
rect 6085 6563 6151 6566
rect 8150 6564 8156 6566
rect 8220 6564 8226 6628
rect 4894 6560 5210 6561
rect 4894 6496 4900 6560
rect 4964 6496 4980 6560
rect 5044 6496 5060 6560
rect 5124 6496 5140 6560
rect 5204 6496 5210 6560
rect 4894 6495 5210 6496
rect 8842 6560 9158 6561
rect 8842 6496 8848 6560
rect 8912 6496 8928 6560
rect 8992 6496 9008 6560
rect 9072 6496 9088 6560
rect 9152 6496 9158 6560
rect 8842 6495 9158 6496
rect 12790 6560 13106 6561
rect 12790 6496 12796 6560
rect 12860 6496 12876 6560
rect 12940 6496 12956 6560
rect 13020 6496 13036 6560
rect 13100 6496 13106 6560
rect 12790 6495 13106 6496
rect 6177 6490 6243 6493
rect 6545 6490 6611 6493
rect 6678 6490 6684 6492
rect 6177 6488 6684 6490
rect 6177 6432 6182 6488
rect 6238 6432 6550 6488
rect 6606 6432 6684 6488
rect 6177 6430 6684 6432
rect 6177 6427 6243 6430
rect 6545 6427 6611 6430
rect 6678 6428 6684 6430
rect 6748 6428 6754 6492
rect 6913 6490 6979 6493
rect 7966 6490 7972 6492
rect 6913 6488 7972 6490
rect 6913 6432 6918 6488
rect 6974 6432 7972 6488
rect 6913 6430 7972 6432
rect 6913 6427 6979 6430
rect 7966 6428 7972 6430
rect 8036 6428 8042 6492
rect 2773 6354 2839 6357
rect 8477 6354 8543 6357
rect 2773 6352 8543 6354
rect 2773 6296 2778 6352
rect 2834 6296 8482 6352
rect 8538 6296 8543 6352
rect 2773 6294 8543 6296
rect 2773 6291 2839 6294
rect 8477 6291 8543 6294
rect 8753 6354 8819 6357
rect 11697 6354 11763 6357
rect 8753 6352 11763 6354
rect 8753 6296 8758 6352
rect 8814 6296 11702 6352
rect 11758 6296 11763 6352
rect 8753 6294 11763 6296
rect 8753 6291 8819 6294
rect 11697 6291 11763 6294
rect 1577 6218 1643 6221
rect 8753 6218 8819 6221
rect 1577 6216 8819 6218
rect 1577 6160 1582 6216
rect 1638 6160 8758 6216
rect 8814 6160 8819 6216
rect 1577 6158 8819 6160
rect 1577 6155 1643 6158
rect 8753 6155 8819 6158
rect 3877 6082 3943 6085
rect 6545 6082 6611 6085
rect 3877 6080 6611 6082
rect 3877 6024 3882 6080
rect 3938 6024 6550 6080
rect 6606 6024 6611 6080
rect 3877 6022 6611 6024
rect 3877 6019 3943 6022
rect 6545 6019 6611 6022
rect 2920 6016 3236 6017
rect 2920 5952 2926 6016
rect 2990 5952 3006 6016
rect 3070 5952 3086 6016
rect 3150 5952 3166 6016
rect 3230 5952 3236 6016
rect 2920 5951 3236 5952
rect 6868 6016 7184 6017
rect 6868 5952 6874 6016
rect 6938 5952 6954 6016
rect 7018 5952 7034 6016
rect 7098 5952 7114 6016
rect 7178 5952 7184 6016
rect 6868 5951 7184 5952
rect 10816 6016 11132 6017
rect 10816 5952 10822 6016
rect 10886 5952 10902 6016
rect 10966 5952 10982 6016
rect 11046 5952 11062 6016
rect 11126 5952 11132 6016
rect 10816 5951 11132 5952
rect 14764 6016 15080 6017
rect 14764 5952 14770 6016
rect 14834 5952 14850 6016
rect 14914 5952 14930 6016
rect 14994 5952 15010 6016
rect 15074 5952 15080 6016
rect 14764 5951 15080 5952
rect 3969 5808 4035 5813
rect 3969 5752 3974 5808
rect 4030 5752 4035 5808
rect 3969 5747 4035 5752
rect 4981 5810 5047 5813
rect 9622 5810 9628 5812
rect 4981 5808 9628 5810
rect 4981 5752 4986 5808
rect 5042 5752 9628 5808
rect 4981 5750 9628 5752
rect 4981 5747 5047 5750
rect 9622 5748 9628 5750
rect 9692 5748 9698 5812
rect 3972 5674 4032 5747
rect 5073 5674 5139 5677
rect 3972 5672 5139 5674
rect 3972 5616 5078 5672
rect 5134 5616 5139 5672
rect 3972 5614 5139 5616
rect 5073 5611 5139 5614
rect 5441 5674 5507 5677
rect 7557 5674 7623 5677
rect 7833 5674 7899 5677
rect 5441 5672 5826 5674
rect 5441 5616 5446 5672
rect 5502 5616 5826 5672
rect 5441 5614 5826 5616
rect 5441 5611 5507 5614
rect 5766 5541 5826 5614
rect 7557 5672 7899 5674
rect 7557 5616 7562 5672
rect 7618 5616 7838 5672
rect 7894 5616 7899 5672
rect 7557 5614 7899 5616
rect 7557 5611 7623 5614
rect 7833 5611 7899 5614
rect 5766 5536 5875 5541
rect 5766 5480 5814 5536
rect 5870 5480 5875 5536
rect 5766 5478 5875 5480
rect 5809 5475 5875 5478
rect 4894 5472 5210 5473
rect 4894 5408 4900 5472
rect 4964 5408 4980 5472
rect 5044 5408 5060 5472
rect 5124 5408 5140 5472
rect 5204 5408 5210 5472
rect 4894 5407 5210 5408
rect 8842 5472 9158 5473
rect 8842 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9008 5472
rect 9072 5408 9088 5472
rect 9152 5408 9158 5472
rect 8842 5407 9158 5408
rect 12790 5472 13106 5473
rect 12790 5408 12796 5472
rect 12860 5408 12876 5472
rect 12940 5408 12956 5472
rect 13020 5408 13036 5472
rect 13100 5408 13106 5472
rect 12790 5407 13106 5408
rect 3049 5402 3115 5405
rect 5349 5404 5415 5405
rect 3550 5402 3556 5404
rect 3049 5400 3556 5402
rect 3049 5344 3054 5400
rect 3110 5344 3556 5400
rect 3049 5342 3556 5344
rect 3049 5339 3115 5342
rect 3550 5340 3556 5342
rect 3620 5340 3626 5404
rect 5349 5402 5396 5404
rect 5304 5400 5396 5402
rect 5304 5344 5354 5400
rect 5304 5342 5396 5344
rect 5349 5340 5396 5342
rect 5460 5340 5466 5404
rect 5625 5402 5691 5405
rect 7649 5402 7715 5405
rect 8477 5404 8543 5405
rect 8477 5402 8524 5404
rect 5625 5400 7715 5402
rect 5625 5344 5630 5400
rect 5686 5344 7654 5400
rect 7710 5344 7715 5400
rect 5625 5342 7715 5344
rect 8432 5400 8524 5402
rect 8432 5344 8482 5400
rect 8432 5342 8524 5344
rect 5349 5339 5415 5340
rect 5625 5339 5691 5342
rect 7649 5339 7715 5342
rect 8477 5340 8524 5342
rect 8588 5340 8594 5404
rect 8477 5339 8543 5340
rect 0 5266 400 5296
rect 3785 5266 3851 5269
rect 0 5264 3851 5266
rect 0 5208 3790 5264
rect 3846 5208 3851 5264
rect 0 5206 3851 5208
rect 0 5176 400 5206
rect 3785 5203 3851 5206
rect 3969 5266 4035 5269
rect 7414 5266 7420 5268
rect 3969 5264 7420 5266
rect 3969 5208 3974 5264
rect 4030 5208 7420 5264
rect 3969 5206 7420 5208
rect 3969 5203 4035 5206
rect 7414 5204 7420 5206
rect 7484 5204 7490 5268
rect 3233 5130 3299 5133
rect 11278 5130 11284 5132
rect 3233 5128 11284 5130
rect 3233 5072 3238 5128
rect 3294 5072 11284 5128
rect 3233 5070 11284 5072
rect 3233 5067 3299 5070
rect 11278 5068 11284 5070
rect 11348 5068 11354 5132
rect 4705 4996 4771 4997
rect 4654 4994 4660 4996
rect 4614 4934 4660 4994
rect 4724 4992 4771 4996
rect 4766 4936 4771 4992
rect 4654 4932 4660 4934
rect 4724 4932 4771 4936
rect 4705 4931 4771 4932
rect 2920 4928 3236 4929
rect 2920 4864 2926 4928
rect 2990 4864 3006 4928
rect 3070 4864 3086 4928
rect 3150 4864 3166 4928
rect 3230 4864 3236 4928
rect 2920 4863 3236 4864
rect 6868 4928 7184 4929
rect 6868 4864 6874 4928
rect 6938 4864 6954 4928
rect 7018 4864 7034 4928
rect 7098 4864 7114 4928
rect 7178 4864 7184 4928
rect 6868 4863 7184 4864
rect 10816 4928 11132 4929
rect 10816 4864 10822 4928
rect 10886 4864 10902 4928
rect 10966 4864 10982 4928
rect 11046 4864 11062 4928
rect 11126 4864 11132 4928
rect 10816 4863 11132 4864
rect 14764 4928 15080 4929
rect 14764 4864 14770 4928
rect 14834 4864 14850 4928
rect 14914 4864 14930 4928
rect 14994 4864 15010 4928
rect 15074 4864 15080 4928
rect 14764 4863 15080 4864
rect 4061 4858 4127 4861
rect 6177 4858 6243 4861
rect 4061 4856 6243 4858
rect 4061 4800 4066 4856
rect 4122 4800 6182 4856
rect 6238 4800 6243 4856
rect 4061 4798 6243 4800
rect 4061 4795 4127 4798
rect 6177 4795 6243 4798
rect 3049 4722 3115 4725
rect 8702 4722 8708 4724
rect 3049 4720 8708 4722
rect 3049 4664 3054 4720
rect 3110 4664 8708 4720
rect 3049 4662 8708 4664
rect 3049 4659 3115 4662
rect 8702 4660 8708 4662
rect 8772 4660 8778 4724
rect 1485 4586 1551 4589
rect 6637 4586 6703 4589
rect 1485 4584 6703 4586
rect 1485 4528 1490 4584
rect 1546 4528 6642 4584
rect 6698 4528 6703 4584
rect 1485 4526 6703 4528
rect 1485 4523 1551 4526
rect 6637 4523 6703 4526
rect 4894 4384 5210 4385
rect 4894 4320 4900 4384
rect 4964 4320 4980 4384
rect 5044 4320 5060 4384
rect 5124 4320 5140 4384
rect 5204 4320 5210 4384
rect 4894 4319 5210 4320
rect 8842 4384 9158 4385
rect 8842 4320 8848 4384
rect 8912 4320 8928 4384
rect 8992 4320 9008 4384
rect 9072 4320 9088 4384
rect 9152 4320 9158 4384
rect 8842 4319 9158 4320
rect 12790 4384 13106 4385
rect 12790 4320 12796 4384
rect 12860 4320 12876 4384
rect 12940 4320 12956 4384
rect 13020 4320 13036 4384
rect 13100 4320 13106 4384
rect 12790 4319 13106 4320
rect 2630 4252 2636 4316
rect 2700 4314 2706 4316
rect 3601 4314 3667 4317
rect 2700 4312 3667 4314
rect 2700 4256 3606 4312
rect 3662 4256 3667 4312
rect 2700 4254 3667 4256
rect 2700 4252 2706 4254
rect 3601 4251 3667 4254
rect 2865 4178 2931 4181
rect 2865 4176 4216 4178
rect 2865 4120 2870 4176
rect 2926 4120 4216 4176
rect 2865 4118 4216 4120
rect 2865 4115 2931 4118
rect 1669 4042 1735 4045
rect 3969 4044 4035 4045
rect 1669 4040 3848 4042
rect 1669 3984 1674 4040
rect 1730 3984 3848 4040
rect 1669 3982 3848 3984
rect 1669 3979 1735 3982
rect 3788 3906 3848 3982
rect 3918 3980 3924 4044
rect 3988 4042 4035 4044
rect 4156 4042 4216 4118
rect 5574 4116 5580 4180
rect 5644 4178 5650 4180
rect 5717 4178 5783 4181
rect 7281 4178 7347 4181
rect 5644 4176 7347 4178
rect 5644 4120 5722 4176
rect 5778 4120 7286 4176
rect 7342 4120 7347 4176
rect 5644 4118 7347 4120
rect 5644 4116 5650 4118
rect 5717 4115 5783 4118
rect 7281 4115 7347 4118
rect 8334 4042 8340 4044
rect 3988 4040 4080 4042
rect 4030 3984 4080 4040
rect 3988 3982 4080 3984
rect 4156 3982 8340 4042
rect 3988 3980 4035 3982
rect 8334 3980 8340 3982
rect 8404 3980 8410 4044
rect 3969 3979 4035 3980
rect 5625 3906 5691 3909
rect 3788 3904 5691 3906
rect 3788 3848 5630 3904
rect 5686 3848 5691 3904
rect 3788 3846 5691 3848
rect 5625 3843 5691 3846
rect 2920 3840 3236 3841
rect 0 3770 400 3800
rect 2920 3776 2926 3840
rect 2990 3776 3006 3840
rect 3070 3776 3086 3840
rect 3150 3776 3166 3840
rect 3230 3776 3236 3840
rect 2920 3775 3236 3776
rect 6868 3840 7184 3841
rect 6868 3776 6874 3840
rect 6938 3776 6954 3840
rect 7018 3776 7034 3840
rect 7098 3776 7114 3840
rect 7178 3776 7184 3840
rect 6868 3775 7184 3776
rect 10816 3840 11132 3841
rect 10816 3776 10822 3840
rect 10886 3776 10902 3840
rect 10966 3776 10982 3840
rect 11046 3776 11062 3840
rect 11126 3776 11132 3840
rect 10816 3775 11132 3776
rect 14764 3840 15080 3841
rect 14764 3776 14770 3840
rect 14834 3776 14850 3840
rect 14914 3776 14930 3840
rect 14994 3776 15010 3840
rect 15074 3776 15080 3840
rect 14764 3775 15080 3776
rect 1393 3770 1459 3773
rect 0 3768 1459 3770
rect 0 3712 1398 3768
rect 1454 3712 1459 3768
rect 0 3710 1459 3712
rect 0 3680 400 3710
rect 1393 3707 1459 3710
rect 2773 3634 2839 3637
rect 4102 3634 4108 3636
rect 2773 3632 4108 3634
rect 2773 3576 2778 3632
rect 2834 3576 4108 3632
rect 2773 3574 4108 3576
rect 2773 3571 2839 3574
rect 4102 3572 4108 3574
rect 4172 3572 4178 3636
rect 2957 3498 3023 3501
rect 3734 3498 3740 3500
rect 2957 3496 3740 3498
rect 2957 3440 2962 3496
rect 3018 3440 3740 3496
rect 2957 3438 3740 3440
rect 2957 3435 3023 3438
rect 3734 3436 3740 3438
rect 3804 3436 3810 3500
rect 1301 3362 1367 3365
rect 3141 3362 3207 3365
rect 1301 3360 3207 3362
rect 1301 3304 1306 3360
rect 1362 3304 3146 3360
rect 3202 3304 3207 3360
rect 1301 3302 3207 3304
rect 1301 3299 1367 3302
rect 3141 3299 3207 3302
rect 4894 3296 5210 3297
rect 4894 3232 4900 3296
rect 4964 3232 4980 3296
rect 5044 3232 5060 3296
rect 5124 3232 5140 3296
rect 5204 3232 5210 3296
rect 4894 3231 5210 3232
rect 8842 3296 9158 3297
rect 8842 3232 8848 3296
rect 8912 3232 8928 3296
rect 8992 3232 9008 3296
rect 9072 3232 9088 3296
rect 9152 3232 9158 3296
rect 8842 3231 9158 3232
rect 12790 3296 13106 3297
rect 12790 3232 12796 3296
rect 12860 3232 12876 3296
rect 12940 3232 12956 3296
rect 13020 3232 13036 3296
rect 13100 3232 13106 3296
rect 12790 3231 13106 3232
rect 2221 3090 2287 3093
rect 9806 3090 9812 3092
rect 2221 3088 9812 3090
rect 2221 3032 2226 3088
rect 2282 3032 9812 3088
rect 2221 3030 9812 3032
rect 2221 3027 2287 3030
rect 9806 3028 9812 3030
rect 9876 3028 9882 3092
rect 2920 2752 3236 2753
rect 2920 2688 2926 2752
rect 2990 2688 3006 2752
rect 3070 2688 3086 2752
rect 3150 2688 3166 2752
rect 3230 2688 3236 2752
rect 2920 2687 3236 2688
rect 6868 2752 7184 2753
rect 6868 2688 6874 2752
rect 6938 2688 6954 2752
rect 7018 2688 7034 2752
rect 7098 2688 7114 2752
rect 7178 2688 7184 2752
rect 6868 2687 7184 2688
rect 10816 2752 11132 2753
rect 10816 2688 10822 2752
rect 10886 2688 10902 2752
rect 10966 2688 10982 2752
rect 11046 2688 11062 2752
rect 11126 2688 11132 2752
rect 10816 2687 11132 2688
rect 14764 2752 15080 2753
rect 14764 2688 14770 2752
rect 14834 2688 14850 2752
rect 14914 2688 14930 2752
rect 14994 2688 15010 2752
rect 15074 2688 15080 2752
rect 14764 2687 15080 2688
rect 0 2274 400 2304
rect 1393 2274 1459 2277
rect 0 2272 1459 2274
rect 0 2216 1398 2272
rect 1454 2216 1459 2272
rect 0 2214 1459 2216
rect 0 2184 400 2214
rect 1393 2211 1459 2214
rect 4894 2208 5210 2209
rect 4894 2144 4900 2208
rect 4964 2144 4980 2208
rect 5044 2144 5060 2208
rect 5124 2144 5140 2208
rect 5204 2144 5210 2208
rect 4894 2143 5210 2144
rect 8842 2208 9158 2209
rect 8842 2144 8848 2208
rect 8912 2144 8928 2208
rect 8992 2144 9008 2208
rect 9072 2144 9088 2208
rect 9152 2144 9158 2208
rect 8842 2143 9158 2144
rect 12790 2208 13106 2209
rect 12790 2144 12796 2208
rect 12860 2144 12876 2208
rect 12940 2144 12956 2208
rect 13020 2144 13036 2208
rect 13100 2144 13106 2208
rect 12790 2143 13106 2144
rect 2920 1664 3236 1665
rect 2920 1600 2926 1664
rect 2990 1600 3006 1664
rect 3070 1600 3086 1664
rect 3150 1600 3166 1664
rect 3230 1600 3236 1664
rect 2920 1599 3236 1600
rect 6868 1664 7184 1665
rect 6868 1600 6874 1664
rect 6938 1600 6954 1664
rect 7018 1600 7034 1664
rect 7098 1600 7114 1664
rect 7178 1600 7184 1664
rect 6868 1599 7184 1600
rect 10816 1664 11132 1665
rect 10816 1600 10822 1664
rect 10886 1600 10902 1664
rect 10966 1600 10982 1664
rect 11046 1600 11062 1664
rect 11126 1600 11132 1664
rect 10816 1599 11132 1600
rect 14764 1664 15080 1665
rect 14764 1600 14770 1664
rect 14834 1600 14850 1664
rect 14914 1600 14930 1664
rect 14994 1600 15010 1664
rect 15074 1600 15080 1664
rect 14764 1599 15080 1600
rect 4894 1120 5210 1121
rect 4894 1056 4900 1120
rect 4964 1056 4980 1120
rect 5044 1056 5060 1120
rect 5124 1056 5140 1120
rect 5204 1056 5210 1120
rect 4894 1055 5210 1056
rect 8842 1120 9158 1121
rect 8842 1056 8848 1120
rect 8912 1056 8928 1120
rect 8992 1056 9008 1120
rect 9072 1056 9088 1120
rect 9152 1056 9158 1120
rect 8842 1055 9158 1056
rect 12790 1120 13106 1121
rect 12790 1056 12796 1120
rect 12860 1056 12876 1120
rect 12940 1056 12956 1120
rect 13020 1056 13036 1120
rect 13100 1056 13106 1120
rect 12790 1055 13106 1056
rect 0 778 400 808
rect 1393 778 1459 781
rect 0 776 1459 778
rect 0 720 1398 776
rect 1454 720 1459 776
rect 0 718 1459 720
rect 0 688 400 718
rect 1393 715 1459 718
<< via3 >>
rect 4900 22876 4964 22880
rect 4900 22820 4904 22876
rect 4904 22820 4960 22876
rect 4960 22820 4964 22876
rect 4900 22816 4964 22820
rect 4980 22876 5044 22880
rect 4980 22820 4984 22876
rect 4984 22820 5040 22876
rect 5040 22820 5044 22876
rect 4980 22816 5044 22820
rect 5060 22876 5124 22880
rect 5060 22820 5064 22876
rect 5064 22820 5120 22876
rect 5120 22820 5124 22876
rect 5060 22816 5124 22820
rect 5140 22876 5204 22880
rect 5140 22820 5144 22876
rect 5144 22820 5200 22876
rect 5200 22820 5204 22876
rect 5140 22816 5204 22820
rect 8848 22876 8912 22880
rect 8848 22820 8852 22876
rect 8852 22820 8908 22876
rect 8908 22820 8912 22876
rect 8848 22816 8912 22820
rect 8928 22876 8992 22880
rect 8928 22820 8932 22876
rect 8932 22820 8988 22876
rect 8988 22820 8992 22876
rect 8928 22816 8992 22820
rect 9008 22876 9072 22880
rect 9008 22820 9012 22876
rect 9012 22820 9068 22876
rect 9068 22820 9072 22876
rect 9008 22816 9072 22820
rect 9088 22876 9152 22880
rect 9088 22820 9092 22876
rect 9092 22820 9148 22876
rect 9148 22820 9152 22876
rect 9088 22816 9152 22820
rect 12796 22876 12860 22880
rect 12796 22820 12800 22876
rect 12800 22820 12856 22876
rect 12856 22820 12860 22876
rect 12796 22816 12860 22820
rect 12876 22876 12940 22880
rect 12876 22820 12880 22876
rect 12880 22820 12936 22876
rect 12936 22820 12940 22876
rect 12876 22816 12940 22820
rect 12956 22876 13020 22880
rect 12956 22820 12960 22876
rect 12960 22820 13016 22876
rect 13016 22820 13020 22876
rect 12956 22816 13020 22820
rect 13036 22876 13100 22880
rect 13036 22820 13040 22876
rect 13040 22820 13096 22876
rect 13096 22820 13100 22876
rect 13036 22816 13100 22820
rect 2926 22332 2990 22336
rect 2926 22276 2930 22332
rect 2930 22276 2986 22332
rect 2986 22276 2990 22332
rect 2926 22272 2990 22276
rect 3006 22332 3070 22336
rect 3006 22276 3010 22332
rect 3010 22276 3066 22332
rect 3066 22276 3070 22332
rect 3006 22272 3070 22276
rect 3086 22332 3150 22336
rect 3086 22276 3090 22332
rect 3090 22276 3146 22332
rect 3146 22276 3150 22332
rect 3086 22272 3150 22276
rect 3166 22332 3230 22336
rect 3166 22276 3170 22332
rect 3170 22276 3226 22332
rect 3226 22276 3230 22332
rect 3166 22272 3230 22276
rect 6874 22332 6938 22336
rect 6874 22276 6878 22332
rect 6878 22276 6934 22332
rect 6934 22276 6938 22332
rect 6874 22272 6938 22276
rect 6954 22332 7018 22336
rect 6954 22276 6958 22332
rect 6958 22276 7014 22332
rect 7014 22276 7018 22332
rect 6954 22272 7018 22276
rect 7034 22332 7098 22336
rect 7034 22276 7038 22332
rect 7038 22276 7094 22332
rect 7094 22276 7098 22332
rect 7034 22272 7098 22276
rect 7114 22332 7178 22336
rect 7114 22276 7118 22332
rect 7118 22276 7174 22332
rect 7174 22276 7178 22332
rect 7114 22272 7178 22276
rect 10822 22332 10886 22336
rect 10822 22276 10826 22332
rect 10826 22276 10882 22332
rect 10882 22276 10886 22332
rect 10822 22272 10886 22276
rect 10902 22332 10966 22336
rect 10902 22276 10906 22332
rect 10906 22276 10962 22332
rect 10962 22276 10966 22332
rect 10902 22272 10966 22276
rect 10982 22332 11046 22336
rect 10982 22276 10986 22332
rect 10986 22276 11042 22332
rect 11042 22276 11046 22332
rect 10982 22272 11046 22276
rect 11062 22332 11126 22336
rect 11062 22276 11066 22332
rect 11066 22276 11122 22332
rect 11122 22276 11126 22332
rect 11062 22272 11126 22276
rect 14770 22332 14834 22336
rect 14770 22276 14774 22332
rect 14774 22276 14830 22332
rect 14830 22276 14834 22332
rect 14770 22272 14834 22276
rect 14850 22332 14914 22336
rect 14850 22276 14854 22332
rect 14854 22276 14910 22332
rect 14910 22276 14914 22332
rect 14850 22272 14914 22276
rect 14930 22332 14994 22336
rect 14930 22276 14934 22332
rect 14934 22276 14990 22332
rect 14990 22276 14994 22332
rect 14930 22272 14994 22276
rect 15010 22332 15074 22336
rect 15010 22276 15014 22332
rect 15014 22276 15070 22332
rect 15070 22276 15074 22332
rect 15010 22272 15074 22276
rect 4900 21788 4964 21792
rect 4900 21732 4904 21788
rect 4904 21732 4960 21788
rect 4960 21732 4964 21788
rect 4900 21728 4964 21732
rect 4980 21788 5044 21792
rect 4980 21732 4984 21788
rect 4984 21732 5040 21788
rect 5040 21732 5044 21788
rect 4980 21728 5044 21732
rect 5060 21788 5124 21792
rect 5060 21732 5064 21788
rect 5064 21732 5120 21788
rect 5120 21732 5124 21788
rect 5060 21728 5124 21732
rect 5140 21788 5204 21792
rect 5140 21732 5144 21788
rect 5144 21732 5200 21788
rect 5200 21732 5204 21788
rect 5140 21728 5204 21732
rect 8848 21788 8912 21792
rect 8848 21732 8852 21788
rect 8852 21732 8908 21788
rect 8908 21732 8912 21788
rect 8848 21728 8912 21732
rect 8928 21788 8992 21792
rect 8928 21732 8932 21788
rect 8932 21732 8988 21788
rect 8988 21732 8992 21788
rect 8928 21728 8992 21732
rect 9008 21788 9072 21792
rect 9008 21732 9012 21788
rect 9012 21732 9068 21788
rect 9068 21732 9072 21788
rect 9008 21728 9072 21732
rect 9088 21788 9152 21792
rect 9088 21732 9092 21788
rect 9092 21732 9148 21788
rect 9148 21732 9152 21788
rect 9088 21728 9152 21732
rect 12796 21788 12860 21792
rect 12796 21732 12800 21788
rect 12800 21732 12856 21788
rect 12856 21732 12860 21788
rect 12796 21728 12860 21732
rect 12876 21788 12940 21792
rect 12876 21732 12880 21788
rect 12880 21732 12936 21788
rect 12936 21732 12940 21788
rect 12876 21728 12940 21732
rect 12956 21788 13020 21792
rect 12956 21732 12960 21788
rect 12960 21732 13016 21788
rect 13016 21732 13020 21788
rect 12956 21728 13020 21732
rect 13036 21788 13100 21792
rect 13036 21732 13040 21788
rect 13040 21732 13096 21788
rect 13096 21732 13100 21788
rect 13036 21728 13100 21732
rect 2926 21244 2990 21248
rect 2926 21188 2930 21244
rect 2930 21188 2986 21244
rect 2986 21188 2990 21244
rect 2926 21184 2990 21188
rect 3006 21244 3070 21248
rect 3006 21188 3010 21244
rect 3010 21188 3066 21244
rect 3066 21188 3070 21244
rect 3006 21184 3070 21188
rect 3086 21244 3150 21248
rect 3086 21188 3090 21244
rect 3090 21188 3146 21244
rect 3146 21188 3150 21244
rect 3086 21184 3150 21188
rect 3166 21244 3230 21248
rect 3166 21188 3170 21244
rect 3170 21188 3226 21244
rect 3226 21188 3230 21244
rect 3166 21184 3230 21188
rect 6874 21244 6938 21248
rect 6874 21188 6878 21244
rect 6878 21188 6934 21244
rect 6934 21188 6938 21244
rect 6874 21184 6938 21188
rect 6954 21244 7018 21248
rect 6954 21188 6958 21244
rect 6958 21188 7014 21244
rect 7014 21188 7018 21244
rect 6954 21184 7018 21188
rect 7034 21244 7098 21248
rect 7034 21188 7038 21244
rect 7038 21188 7094 21244
rect 7094 21188 7098 21244
rect 7034 21184 7098 21188
rect 7114 21244 7178 21248
rect 7114 21188 7118 21244
rect 7118 21188 7174 21244
rect 7174 21188 7178 21244
rect 7114 21184 7178 21188
rect 10822 21244 10886 21248
rect 10822 21188 10826 21244
rect 10826 21188 10882 21244
rect 10882 21188 10886 21244
rect 10822 21184 10886 21188
rect 10902 21244 10966 21248
rect 10902 21188 10906 21244
rect 10906 21188 10962 21244
rect 10962 21188 10966 21244
rect 10902 21184 10966 21188
rect 10982 21244 11046 21248
rect 10982 21188 10986 21244
rect 10986 21188 11042 21244
rect 11042 21188 11046 21244
rect 10982 21184 11046 21188
rect 11062 21244 11126 21248
rect 11062 21188 11066 21244
rect 11066 21188 11122 21244
rect 11122 21188 11126 21244
rect 11062 21184 11126 21188
rect 14770 21244 14834 21248
rect 14770 21188 14774 21244
rect 14774 21188 14830 21244
rect 14830 21188 14834 21244
rect 14770 21184 14834 21188
rect 14850 21244 14914 21248
rect 14850 21188 14854 21244
rect 14854 21188 14910 21244
rect 14910 21188 14914 21244
rect 14850 21184 14914 21188
rect 14930 21244 14994 21248
rect 14930 21188 14934 21244
rect 14934 21188 14990 21244
rect 14990 21188 14994 21244
rect 14930 21184 14994 21188
rect 15010 21244 15074 21248
rect 15010 21188 15014 21244
rect 15014 21188 15070 21244
rect 15070 21188 15074 21244
rect 15010 21184 15074 21188
rect 4900 20700 4964 20704
rect 4900 20644 4904 20700
rect 4904 20644 4960 20700
rect 4960 20644 4964 20700
rect 4900 20640 4964 20644
rect 4980 20700 5044 20704
rect 4980 20644 4984 20700
rect 4984 20644 5040 20700
rect 5040 20644 5044 20700
rect 4980 20640 5044 20644
rect 5060 20700 5124 20704
rect 5060 20644 5064 20700
rect 5064 20644 5120 20700
rect 5120 20644 5124 20700
rect 5060 20640 5124 20644
rect 5140 20700 5204 20704
rect 5140 20644 5144 20700
rect 5144 20644 5200 20700
rect 5200 20644 5204 20700
rect 5140 20640 5204 20644
rect 8848 20700 8912 20704
rect 8848 20644 8852 20700
rect 8852 20644 8908 20700
rect 8908 20644 8912 20700
rect 8848 20640 8912 20644
rect 8928 20700 8992 20704
rect 8928 20644 8932 20700
rect 8932 20644 8988 20700
rect 8988 20644 8992 20700
rect 8928 20640 8992 20644
rect 9008 20700 9072 20704
rect 9008 20644 9012 20700
rect 9012 20644 9068 20700
rect 9068 20644 9072 20700
rect 9008 20640 9072 20644
rect 9088 20700 9152 20704
rect 9088 20644 9092 20700
rect 9092 20644 9148 20700
rect 9148 20644 9152 20700
rect 9088 20640 9152 20644
rect 12796 20700 12860 20704
rect 12796 20644 12800 20700
rect 12800 20644 12856 20700
rect 12856 20644 12860 20700
rect 12796 20640 12860 20644
rect 12876 20700 12940 20704
rect 12876 20644 12880 20700
rect 12880 20644 12936 20700
rect 12936 20644 12940 20700
rect 12876 20640 12940 20644
rect 12956 20700 13020 20704
rect 12956 20644 12960 20700
rect 12960 20644 13016 20700
rect 13016 20644 13020 20700
rect 12956 20640 13020 20644
rect 13036 20700 13100 20704
rect 13036 20644 13040 20700
rect 13040 20644 13096 20700
rect 13096 20644 13100 20700
rect 13036 20640 13100 20644
rect 2926 20156 2990 20160
rect 2926 20100 2930 20156
rect 2930 20100 2986 20156
rect 2986 20100 2990 20156
rect 2926 20096 2990 20100
rect 3006 20156 3070 20160
rect 3006 20100 3010 20156
rect 3010 20100 3066 20156
rect 3066 20100 3070 20156
rect 3006 20096 3070 20100
rect 3086 20156 3150 20160
rect 3086 20100 3090 20156
rect 3090 20100 3146 20156
rect 3146 20100 3150 20156
rect 3086 20096 3150 20100
rect 3166 20156 3230 20160
rect 3166 20100 3170 20156
rect 3170 20100 3226 20156
rect 3226 20100 3230 20156
rect 3166 20096 3230 20100
rect 6874 20156 6938 20160
rect 6874 20100 6878 20156
rect 6878 20100 6934 20156
rect 6934 20100 6938 20156
rect 6874 20096 6938 20100
rect 6954 20156 7018 20160
rect 6954 20100 6958 20156
rect 6958 20100 7014 20156
rect 7014 20100 7018 20156
rect 6954 20096 7018 20100
rect 7034 20156 7098 20160
rect 7034 20100 7038 20156
rect 7038 20100 7094 20156
rect 7094 20100 7098 20156
rect 7034 20096 7098 20100
rect 7114 20156 7178 20160
rect 7114 20100 7118 20156
rect 7118 20100 7174 20156
rect 7174 20100 7178 20156
rect 7114 20096 7178 20100
rect 10822 20156 10886 20160
rect 10822 20100 10826 20156
rect 10826 20100 10882 20156
rect 10882 20100 10886 20156
rect 10822 20096 10886 20100
rect 10902 20156 10966 20160
rect 10902 20100 10906 20156
rect 10906 20100 10962 20156
rect 10962 20100 10966 20156
rect 10902 20096 10966 20100
rect 10982 20156 11046 20160
rect 10982 20100 10986 20156
rect 10986 20100 11042 20156
rect 11042 20100 11046 20156
rect 10982 20096 11046 20100
rect 11062 20156 11126 20160
rect 11062 20100 11066 20156
rect 11066 20100 11122 20156
rect 11122 20100 11126 20156
rect 11062 20096 11126 20100
rect 14770 20156 14834 20160
rect 14770 20100 14774 20156
rect 14774 20100 14830 20156
rect 14830 20100 14834 20156
rect 14770 20096 14834 20100
rect 14850 20156 14914 20160
rect 14850 20100 14854 20156
rect 14854 20100 14910 20156
rect 14910 20100 14914 20156
rect 14850 20096 14914 20100
rect 14930 20156 14994 20160
rect 14930 20100 14934 20156
rect 14934 20100 14990 20156
rect 14990 20100 14994 20156
rect 14930 20096 14994 20100
rect 15010 20156 15074 20160
rect 15010 20100 15014 20156
rect 15014 20100 15070 20156
rect 15070 20100 15074 20156
rect 15010 20096 15074 20100
rect 4900 19612 4964 19616
rect 4900 19556 4904 19612
rect 4904 19556 4960 19612
rect 4960 19556 4964 19612
rect 4900 19552 4964 19556
rect 4980 19612 5044 19616
rect 4980 19556 4984 19612
rect 4984 19556 5040 19612
rect 5040 19556 5044 19612
rect 4980 19552 5044 19556
rect 5060 19612 5124 19616
rect 5060 19556 5064 19612
rect 5064 19556 5120 19612
rect 5120 19556 5124 19612
rect 5060 19552 5124 19556
rect 5140 19612 5204 19616
rect 5140 19556 5144 19612
rect 5144 19556 5200 19612
rect 5200 19556 5204 19612
rect 5140 19552 5204 19556
rect 8848 19612 8912 19616
rect 8848 19556 8852 19612
rect 8852 19556 8908 19612
rect 8908 19556 8912 19612
rect 8848 19552 8912 19556
rect 8928 19612 8992 19616
rect 8928 19556 8932 19612
rect 8932 19556 8988 19612
rect 8988 19556 8992 19612
rect 8928 19552 8992 19556
rect 9008 19612 9072 19616
rect 9008 19556 9012 19612
rect 9012 19556 9068 19612
rect 9068 19556 9072 19612
rect 9008 19552 9072 19556
rect 9088 19612 9152 19616
rect 9088 19556 9092 19612
rect 9092 19556 9148 19612
rect 9148 19556 9152 19612
rect 9088 19552 9152 19556
rect 12796 19612 12860 19616
rect 12796 19556 12800 19612
rect 12800 19556 12856 19612
rect 12856 19556 12860 19612
rect 12796 19552 12860 19556
rect 12876 19612 12940 19616
rect 12876 19556 12880 19612
rect 12880 19556 12936 19612
rect 12936 19556 12940 19612
rect 12876 19552 12940 19556
rect 12956 19612 13020 19616
rect 12956 19556 12960 19612
rect 12960 19556 13016 19612
rect 13016 19556 13020 19612
rect 12956 19552 13020 19556
rect 13036 19612 13100 19616
rect 13036 19556 13040 19612
rect 13040 19556 13096 19612
rect 13096 19556 13100 19612
rect 13036 19552 13100 19556
rect 2926 19068 2990 19072
rect 2926 19012 2930 19068
rect 2930 19012 2986 19068
rect 2986 19012 2990 19068
rect 2926 19008 2990 19012
rect 3006 19068 3070 19072
rect 3006 19012 3010 19068
rect 3010 19012 3066 19068
rect 3066 19012 3070 19068
rect 3006 19008 3070 19012
rect 3086 19068 3150 19072
rect 3086 19012 3090 19068
rect 3090 19012 3146 19068
rect 3146 19012 3150 19068
rect 3086 19008 3150 19012
rect 3166 19068 3230 19072
rect 3166 19012 3170 19068
rect 3170 19012 3226 19068
rect 3226 19012 3230 19068
rect 3166 19008 3230 19012
rect 6874 19068 6938 19072
rect 6874 19012 6878 19068
rect 6878 19012 6934 19068
rect 6934 19012 6938 19068
rect 6874 19008 6938 19012
rect 6954 19068 7018 19072
rect 6954 19012 6958 19068
rect 6958 19012 7014 19068
rect 7014 19012 7018 19068
rect 6954 19008 7018 19012
rect 7034 19068 7098 19072
rect 7034 19012 7038 19068
rect 7038 19012 7094 19068
rect 7094 19012 7098 19068
rect 7034 19008 7098 19012
rect 7114 19068 7178 19072
rect 7114 19012 7118 19068
rect 7118 19012 7174 19068
rect 7174 19012 7178 19068
rect 7114 19008 7178 19012
rect 10822 19068 10886 19072
rect 10822 19012 10826 19068
rect 10826 19012 10882 19068
rect 10882 19012 10886 19068
rect 10822 19008 10886 19012
rect 10902 19068 10966 19072
rect 10902 19012 10906 19068
rect 10906 19012 10962 19068
rect 10962 19012 10966 19068
rect 10902 19008 10966 19012
rect 10982 19068 11046 19072
rect 10982 19012 10986 19068
rect 10986 19012 11042 19068
rect 11042 19012 11046 19068
rect 10982 19008 11046 19012
rect 11062 19068 11126 19072
rect 11062 19012 11066 19068
rect 11066 19012 11122 19068
rect 11122 19012 11126 19068
rect 11062 19008 11126 19012
rect 14770 19068 14834 19072
rect 14770 19012 14774 19068
rect 14774 19012 14830 19068
rect 14830 19012 14834 19068
rect 14770 19008 14834 19012
rect 14850 19068 14914 19072
rect 14850 19012 14854 19068
rect 14854 19012 14910 19068
rect 14910 19012 14914 19068
rect 14850 19008 14914 19012
rect 14930 19068 14994 19072
rect 14930 19012 14934 19068
rect 14934 19012 14990 19068
rect 14990 19012 14994 19068
rect 14930 19008 14994 19012
rect 15010 19068 15074 19072
rect 15010 19012 15014 19068
rect 15014 19012 15070 19068
rect 15070 19012 15074 19068
rect 15010 19008 15074 19012
rect 4900 18524 4964 18528
rect 4900 18468 4904 18524
rect 4904 18468 4960 18524
rect 4960 18468 4964 18524
rect 4900 18464 4964 18468
rect 4980 18524 5044 18528
rect 4980 18468 4984 18524
rect 4984 18468 5040 18524
rect 5040 18468 5044 18524
rect 4980 18464 5044 18468
rect 5060 18524 5124 18528
rect 5060 18468 5064 18524
rect 5064 18468 5120 18524
rect 5120 18468 5124 18524
rect 5060 18464 5124 18468
rect 5140 18524 5204 18528
rect 5140 18468 5144 18524
rect 5144 18468 5200 18524
rect 5200 18468 5204 18524
rect 5140 18464 5204 18468
rect 8848 18524 8912 18528
rect 8848 18468 8852 18524
rect 8852 18468 8908 18524
rect 8908 18468 8912 18524
rect 8848 18464 8912 18468
rect 8928 18524 8992 18528
rect 8928 18468 8932 18524
rect 8932 18468 8988 18524
rect 8988 18468 8992 18524
rect 8928 18464 8992 18468
rect 9008 18524 9072 18528
rect 9008 18468 9012 18524
rect 9012 18468 9068 18524
rect 9068 18468 9072 18524
rect 9008 18464 9072 18468
rect 9088 18524 9152 18528
rect 9088 18468 9092 18524
rect 9092 18468 9148 18524
rect 9148 18468 9152 18524
rect 9088 18464 9152 18468
rect 12796 18524 12860 18528
rect 12796 18468 12800 18524
rect 12800 18468 12856 18524
rect 12856 18468 12860 18524
rect 12796 18464 12860 18468
rect 12876 18524 12940 18528
rect 12876 18468 12880 18524
rect 12880 18468 12936 18524
rect 12936 18468 12940 18524
rect 12876 18464 12940 18468
rect 12956 18524 13020 18528
rect 12956 18468 12960 18524
rect 12960 18468 13016 18524
rect 13016 18468 13020 18524
rect 12956 18464 13020 18468
rect 13036 18524 13100 18528
rect 13036 18468 13040 18524
rect 13040 18468 13096 18524
rect 13096 18468 13100 18524
rect 13036 18464 13100 18468
rect 2926 17980 2990 17984
rect 2926 17924 2930 17980
rect 2930 17924 2986 17980
rect 2986 17924 2990 17980
rect 2926 17920 2990 17924
rect 3006 17980 3070 17984
rect 3006 17924 3010 17980
rect 3010 17924 3066 17980
rect 3066 17924 3070 17980
rect 3006 17920 3070 17924
rect 3086 17980 3150 17984
rect 3086 17924 3090 17980
rect 3090 17924 3146 17980
rect 3146 17924 3150 17980
rect 3086 17920 3150 17924
rect 3166 17980 3230 17984
rect 3166 17924 3170 17980
rect 3170 17924 3226 17980
rect 3226 17924 3230 17980
rect 3166 17920 3230 17924
rect 6874 17980 6938 17984
rect 6874 17924 6878 17980
rect 6878 17924 6934 17980
rect 6934 17924 6938 17980
rect 6874 17920 6938 17924
rect 6954 17980 7018 17984
rect 6954 17924 6958 17980
rect 6958 17924 7014 17980
rect 7014 17924 7018 17980
rect 6954 17920 7018 17924
rect 7034 17980 7098 17984
rect 7034 17924 7038 17980
rect 7038 17924 7094 17980
rect 7094 17924 7098 17980
rect 7034 17920 7098 17924
rect 7114 17980 7178 17984
rect 7114 17924 7118 17980
rect 7118 17924 7174 17980
rect 7174 17924 7178 17980
rect 7114 17920 7178 17924
rect 10822 17980 10886 17984
rect 10822 17924 10826 17980
rect 10826 17924 10882 17980
rect 10882 17924 10886 17980
rect 10822 17920 10886 17924
rect 10902 17980 10966 17984
rect 10902 17924 10906 17980
rect 10906 17924 10962 17980
rect 10962 17924 10966 17980
rect 10902 17920 10966 17924
rect 10982 17980 11046 17984
rect 10982 17924 10986 17980
rect 10986 17924 11042 17980
rect 11042 17924 11046 17980
rect 10982 17920 11046 17924
rect 11062 17980 11126 17984
rect 11062 17924 11066 17980
rect 11066 17924 11122 17980
rect 11122 17924 11126 17980
rect 11062 17920 11126 17924
rect 14770 17980 14834 17984
rect 14770 17924 14774 17980
rect 14774 17924 14830 17980
rect 14830 17924 14834 17980
rect 14770 17920 14834 17924
rect 14850 17980 14914 17984
rect 14850 17924 14854 17980
rect 14854 17924 14910 17980
rect 14910 17924 14914 17980
rect 14850 17920 14914 17924
rect 14930 17980 14994 17984
rect 14930 17924 14934 17980
rect 14934 17924 14990 17980
rect 14990 17924 14994 17980
rect 14930 17920 14994 17924
rect 15010 17980 15074 17984
rect 15010 17924 15014 17980
rect 15014 17924 15070 17980
rect 15070 17924 15074 17980
rect 15010 17920 15074 17924
rect 4900 17436 4964 17440
rect 4900 17380 4904 17436
rect 4904 17380 4960 17436
rect 4960 17380 4964 17436
rect 4900 17376 4964 17380
rect 4980 17436 5044 17440
rect 4980 17380 4984 17436
rect 4984 17380 5040 17436
rect 5040 17380 5044 17436
rect 4980 17376 5044 17380
rect 5060 17436 5124 17440
rect 5060 17380 5064 17436
rect 5064 17380 5120 17436
rect 5120 17380 5124 17436
rect 5060 17376 5124 17380
rect 5140 17436 5204 17440
rect 5140 17380 5144 17436
rect 5144 17380 5200 17436
rect 5200 17380 5204 17436
rect 5140 17376 5204 17380
rect 8848 17436 8912 17440
rect 8848 17380 8852 17436
rect 8852 17380 8908 17436
rect 8908 17380 8912 17436
rect 8848 17376 8912 17380
rect 8928 17436 8992 17440
rect 8928 17380 8932 17436
rect 8932 17380 8988 17436
rect 8988 17380 8992 17436
rect 8928 17376 8992 17380
rect 9008 17436 9072 17440
rect 9008 17380 9012 17436
rect 9012 17380 9068 17436
rect 9068 17380 9072 17436
rect 9008 17376 9072 17380
rect 9088 17436 9152 17440
rect 9088 17380 9092 17436
rect 9092 17380 9148 17436
rect 9148 17380 9152 17436
rect 9088 17376 9152 17380
rect 12796 17436 12860 17440
rect 12796 17380 12800 17436
rect 12800 17380 12856 17436
rect 12856 17380 12860 17436
rect 12796 17376 12860 17380
rect 12876 17436 12940 17440
rect 12876 17380 12880 17436
rect 12880 17380 12936 17436
rect 12936 17380 12940 17436
rect 12876 17376 12940 17380
rect 12956 17436 13020 17440
rect 12956 17380 12960 17436
rect 12960 17380 13016 17436
rect 13016 17380 13020 17436
rect 12956 17376 13020 17380
rect 13036 17436 13100 17440
rect 13036 17380 13040 17436
rect 13040 17380 13096 17436
rect 13096 17380 13100 17436
rect 13036 17376 13100 17380
rect 2926 16892 2990 16896
rect 2926 16836 2930 16892
rect 2930 16836 2986 16892
rect 2986 16836 2990 16892
rect 2926 16832 2990 16836
rect 3006 16892 3070 16896
rect 3006 16836 3010 16892
rect 3010 16836 3066 16892
rect 3066 16836 3070 16892
rect 3006 16832 3070 16836
rect 3086 16892 3150 16896
rect 3086 16836 3090 16892
rect 3090 16836 3146 16892
rect 3146 16836 3150 16892
rect 3086 16832 3150 16836
rect 3166 16892 3230 16896
rect 3166 16836 3170 16892
rect 3170 16836 3226 16892
rect 3226 16836 3230 16892
rect 3166 16832 3230 16836
rect 6874 16892 6938 16896
rect 6874 16836 6878 16892
rect 6878 16836 6934 16892
rect 6934 16836 6938 16892
rect 6874 16832 6938 16836
rect 6954 16892 7018 16896
rect 6954 16836 6958 16892
rect 6958 16836 7014 16892
rect 7014 16836 7018 16892
rect 6954 16832 7018 16836
rect 7034 16892 7098 16896
rect 7034 16836 7038 16892
rect 7038 16836 7094 16892
rect 7094 16836 7098 16892
rect 7034 16832 7098 16836
rect 7114 16892 7178 16896
rect 7114 16836 7118 16892
rect 7118 16836 7174 16892
rect 7174 16836 7178 16892
rect 7114 16832 7178 16836
rect 10822 16892 10886 16896
rect 10822 16836 10826 16892
rect 10826 16836 10882 16892
rect 10882 16836 10886 16892
rect 10822 16832 10886 16836
rect 10902 16892 10966 16896
rect 10902 16836 10906 16892
rect 10906 16836 10962 16892
rect 10962 16836 10966 16892
rect 10902 16832 10966 16836
rect 10982 16892 11046 16896
rect 10982 16836 10986 16892
rect 10986 16836 11042 16892
rect 11042 16836 11046 16892
rect 10982 16832 11046 16836
rect 11062 16892 11126 16896
rect 11062 16836 11066 16892
rect 11066 16836 11122 16892
rect 11122 16836 11126 16892
rect 11062 16832 11126 16836
rect 14770 16892 14834 16896
rect 14770 16836 14774 16892
rect 14774 16836 14830 16892
rect 14830 16836 14834 16892
rect 14770 16832 14834 16836
rect 14850 16892 14914 16896
rect 14850 16836 14854 16892
rect 14854 16836 14910 16892
rect 14910 16836 14914 16892
rect 14850 16832 14914 16836
rect 14930 16892 14994 16896
rect 14930 16836 14934 16892
rect 14934 16836 14990 16892
rect 14990 16836 14994 16892
rect 14930 16832 14994 16836
rect 15010 16892 15074 16896
rect 15010 16836 15014 16892
rect 15014 16836 15070 16892
rect 15070 16836 15074 16892
rect 15010 16832 15074 16836
rect 4900 16348 4964 16352
rect 4900 16292 4904 16348
rect 4904 16292 4960 16348
rect 4960 16292 4964 16348
rect 4900 16288 4964 16292
rect 4980 16348 5044 16352
rect 4980 16292 4984 16348
rect 4984 16292 5040 16348
rect 5040 16292 5044 16348
rect 4980 16288 5044 16292
rect 5060 16348 5124 16352
rect 5060 16292 5064 16348
rect 5064 16292 5120 16348
rect 5120 16292 5124 16348
rect 5060 16288 5124 16292
rect 5140 16348 5204 16352
rect 5140 16292 5144 16348
rect 5144 16292 5200 16348
rect 5200 16292 5204 16348
rect 5140 16288 5204 16292
rect 8848 16348 8912 16352
rect 8848 16292 8852 16348
rect 8852 16292 8908 16348
rect 8908 16292 8912 16348
rect 8848 16288 8912 16292
rect 8928 16348 8992 16352
rect 8928 16292 8932 16348
rect 8932 16292 8988 16348
rect 8988 16292 8992 16348
rect 8928 16288 8992 16292
rect 9008 16348 9072 16352
rect 9008 16292 9012 16348
rect 9012 16292 9068 16348
rect 9068 16292 9072 16348
rect 9008 16288 9072 16292
rect 9088 16348 9152 16352
rect 9088 16292 9092 16348
rect 9092 16292 9148 16348
rect 9148 16292 9152 16348
rect 9088 16288 9152 16292
rect 12796 16348 12860 16352
rect 12796 16292 12800 16348
rect 12800 16292 12856 16348
rect 12856 16292 12860 16348
rect 12796 16288 12860 16292
rect 12876 16348 12940 16352
rect 12876 16292 12880 16348
rect 12880 16292 12936 16348
rect 12936 16292 12940 16348
rect 12876 16288 12940 16292
rect 12956 16348 13020 16352
rect 12956 16292 12960 16348
rect 12960 16292 13016 16348
rect 13016 16292 13020 16348
rect 12956 16288 13020 16292
rect 13036 16348 13100 16352
rect 13036 16292 13040 16348
rect 13040 16292 13096 16348
rect 13096 16292 13100 16348
rect 13036 16288 13100 16292
rect 2926 15804 2990 15808
rect 2926 15748 2930 15804
rect 2930 15748 2986 15804
rect 2986 15748 2990 15804
rect 2926 15744 2990 15748
rect 3006 15804 3070 15808
rect 3006 15748 3010 15804
rect 3010 15748 3066 15804
rect 3066 15748 3070 15804
rect 3006 15744 3070 15748
rect 3086 15804 3150 15808
rect 3086 15748 3090 15804
rect 3090 15748 3146 15804
rect 3146 15748 3150 15804
rect 3086 15744 3150 15748
rect 3166 15804 3230 15808
rect 3166 15748 3170 15804
rect 3170 15748 3226 15804
rect 3226 15748 3230 15804
rect 3166 15744 3230 15748
rect 6874 15804 6938 15808
rect 6874 15748 6878 15804
rect 6878 15748 6934 15804
rect 6934 15748 6938 15804
rect 6874 15744 6938 15748
rect 6954 15804 7018 15808
rect 6954 15748 6958 15804
rect 6958 15748 7014 15804
rect 7014 15748 7018 15804
rect 6954 15744 7018 15748
rect 7034 15804 7098 15808
rect 7034 15748 7038 15804
rect 7038 15748 7094 15804
rect 7094 15748 7098 15804
rect 7034 15744 7098 15748
rect 7114 15804 7178 15808
rect 7114 15748 7118 15804
rect 7118 15748 7174 15804
rect 7174 15748 7178 15804
rect 7114 15744 7178 15748
rect 10822 15804 10886 15808
rect 10822 15748 10826 15804
rect 10826 15748 10882 15804
rect 10882 15748 10886 15804
rect 10822 15744 10886 15748
rect 10902 15804 10966 15808
rect 10902 15748 10906 15804
rect 10906 15748 10962 15804
rect 10962 15748 10966 15804
rect 10902 15744 10966 15748
rect 10982 15804 11046 15808
rect 10982 15748 10986 15804
rect 10986 15748 11042 15804
rect 11042 15748 11046 15804
rect 10982 15744 11046 15748
rect 11062 15804 11126 15808
rect 11062 15748 11066 15804
rect 11066 15748 11122 15804
rect 11122 15748 11126 15804
rect 11062 15744 11126 15748
rect 14770 15804 14834 15808
rect 14770 15748 14774 15804
rect 14774 15748 14830 15804
rect 14830 15748 14834 15804
rect 14770 15744 14834 15748
rect 14850 15804 14914 15808
rect 14850 15748 14854 15804
rect 14854 15748 14910 15804
rect 14910 15748 14914 15804
rect 14850 15744 14914 15748
rect 14930 15804 14994 15808
rect 14930 15748 14934 15804
rect 14934 15748 14990 15804
rect 14990 15748 14994 15804
rect 14930 15744 14994 15748
rect 15010 15804 15074 15808
rect 15010 15748 15014 15804
rect 15014 15748 15070 15804
rect 15070 15748 15074 15804
rect 15010 15744 15074 15748
rect 5396 15404 5460 15468
rect 6500 15404 6564 15468
rect 4900 15260 4964 15264
rect 4900 15204 4904 15260
rect 4904 15204 4960 15260
rect 4960 15204 4964 15260
rect 4900 15200 4964 15204
rect 4980 15260 5044 15264
rect 4980 15204 4984 15260
rect 4984 15204 5040 15260
rect 5040 15204 5044 15260
rect 4980 15200 5044 15204
rect 5060 15260 5124 15264
rect 5060 15204 5064 15260
rect 5064 15204 5120 15260
rect 5120 15204 5124 15260
rect 5060 15200 5124 15204
rect 5140 15260 5204 15264
rect 5140 15204 5144 15260
rect 5144 15204 5200 15260
rect 5200 15204 5204 15260
rect 5140 15200 5204 15204
rect 8848 15260 8912 15264
rect 8848 15204 8852 15260
rect 8852 15204 8908 15260
rect 8908 15204 8912 15260
rect 8848 15200 8912 15204
rect 8928 15260 8992 15264
rect 8928 15204 8932 15260
rect 8932 15204 8988 15260
rect 8988 15204 8992 15260
rect 8928 15200 8992 15204
rect 9008 15260 9072 15264
rect 9008 15204 9012 15260
rect 9012 15204 9068 15260
rect 9068 15204 9072 15260
rect 9008 15200 9072 15204
rect 9088 15260 9152 15264
rect 9088 15204 9092 15260
rect 9092 15204 9148 15260
rect 9148 15204 9152 15260
rect 9088 15200 9152 15204
rect 12796 15260 12860 15264
rect 12796 15204 12800 15260
rect 12800 15204 12856 15260
rect 12856 15204 12860 15260
rect 12796 15200 12860 15204
rect 12876 15260 12940 15264
rect 12876 15204 12880 15260
rect 12880 15204 12936 15260
rect 12936 15204 12940 15260
rect 12876 15200 12940 15204
rect 12956 15260 13020 15264
rect 12956 15204 12960 15260
rect 12960 15204 13016 15260
rect 13016 15204 13020 15260
rect 12956 15200 13020 15204
rect 13036 15260 13100 15264
rect 13036 15204 13040 15260
rect 13040 15204 13096 15260
rect 13096 15204 13100 15260
rect 13036 15200 13100 15204
rect 7420 14860 7484 14924
rect 2926 14716 2990 14720
rect 2926 14660 2930 14716
rect 2930 14660 2986 14716
rect 2986 14660 2990 14716
rect 2926 14656 2990 14660
rect 3006 14716 3070 14720
rect 3006 14660 3010 14716
rect 3010 14660 3066 14716
rect 3066 14660 3070 14716
rect 3006 14656 3070 14660
rect 3086 14716 3150 14720
rect 3086 14660 3090 14716
rect 3090 14660 3146 14716
rect 3146 14660 3150 14716
rect 3086 14656 3150 14660
rect 3166 14716 3230 14720
rect 3166 14660 3170 14716
rect 3170 14660 3226 14716
rect 3226 14660 3230 14716
rect 3166 14656 3230 14660
rect 6874 14716 6938 14720
rect 6874 14660 6878 14716
rect 6878 14660 6934 14716
rect 6934 14660 6938 14716
rect 6874 14656 6938 14660
rect 6954 14716 7018 14720
rect 6954 14660 6958 14716
rect 6958 14660 7014 14716
rect 7014 14660 7018 14716
rect 6954 14656 7018 14660
rect 7034 14716 7098 14720
rect 7034 14660 7038 14716
rect 7038 14660 7094 14716
rect 7094 14660 7098 14716
rect 7034 14656 7098 14660
rect 7114 14716 7178 14720
rect 7114 14660 7118 14716
rect 7118 14660 7174 14716
rect 7174 14660 7178 14716
rect 7114 14656 7178 14660
rect 10822 14716 10886 14720
rect 10822 14660 10826 14716
rect 10826 14660 10882 14716
rect 10882 14660 10886 14716
rect 10822 14656 10886 14660
rect 10902 14716 10966 14720
rect 10902 14660 10906 14716
rect 10906 14660 10962 14716
rect 10962 14660 10966 14716
rect 10902 14656 10966 14660
rect 10982 14716 11046 14720
rect 10982 14660 10986 14716
rect 10986 14660 11042 14716
rect 11042 14660 11046 14716
rect 10982 14656 11046 14660
rect 11062 14716 11126 14720
rect 11062 14660 11066 14716
rect 11066 14660 11122 14716
rect 11122 14660 11126 14716
rect 11062 14656 11126 14660
rect 14770 14716 14834 14720
rect 14770 14660 14774 14716
rect 14774 14660 14830 14716
rect 14830 14660 14834 14716
rect 14770 14656 14834 14660
rect 14850 14716 14914 14720
rect 14850 14660 14854 14716
rect 14854 14660 14910 14716
rect 14910 14660 14914 14716
rect 14850 14656 14914 14660
rect 14930 14716 14994 14720
rect 14930 14660 14934 14716
rect 14934 14660 14990 14716
rect 14990 14660 14994 14716
rect 14930 14656 14994 14660
rect 15010 14716 15074 14720
rect 15010 14660 15014 14716
rect 15014 14660 15070 14716
rect 15070 14660 15074 14716
rect 15010 14656 15074 14660
rect 3924 14316 3988 14380
rect 4900 14172 4964 14176
rect 4900 14116 4904 14172
rect 4904 14116 4960 14172
rect 4960 14116 4964 14172
rect 4900 14112 4964 14116
rect 4980 14172 5044 14176
rect 4980 14116 4984 14172
rect 4984 14116 5040 14172
rect 5040 14116 5044 14172
rect 4980 14112 5044 14116
rect 5060 14172 5124 14176
rect 5060 14116 5064 14172
rect 5064 14116 5120 14172
rect 5120 14116 5124 14172
rect 5060 14112 5124 14116
rect 5140 14172 5204 14176
rect 5140 14116 5144 14172
rect 5144 14116 5200 14172
rect 5200 14116 5204 14172
rect 5140 14112 5204 14116
rect 8848 14172 8912 14176
rect 8848 14116 8852 14172
rect 8852 14116 8908 14172
rect 8908 14116 8912 14172
rect 8848 14112 8912 14116
rect 8928 14172 8992 14176
rect 8928 14116 8932 14172
rect 8932 14116 8988 14172
rect 8988 14116 8992 14172
rect 8928 14112 8992 14116
rect 9008 14172 9072 14176
rect 9008 14116 9012 14172
rect 9012 14116 9068 14172
rect 9068 14116 9072 14172
rect 9008 14112 9072 14116
rect 9088 14172 9152 14176
rect 9088 14116 9092 14172
rect 9092 14116 9148 14172
rect 9148 14116 9152 14172
rect 9088 14112 9152 14116
rect 12796 14172 12860 14176
rect 12796 14116 12800 14172
rect 12800 14116 12856 14172
rect 12856 14116 12860 14172
rect 12796 14112 12860 14116
rect 12876 14172 12940 14176
rect 12876 14116 12880 14172
rect 12880 14116 12936 14172
rect 12936 14116 12940 14172
rect 12876 14112 12940 14116
rect 12956 14172 13020 14176
rect 12956 14116 12960 14172
rect 12960 14116 13016 14172
rect 13016 14116 13020 14172
rect 12956 14112 13020 14116
rect 13036 14172 13100 14176
rect 13036 14116 13040 14172
rect 13040 14116 13096 14172
rect 13096 14116 13100 14172
rect 13036 14112 13100 14116
rect 2926 13628 2990 13632
rect 2926 13572 2930 13628
rect 2930 13572 2986 13628
rect 2986 13572 2990 13628
rect 2926 13568 2990 13572
rect 3006 13628 3070 13632
rect 3006 13572 3010 13628
rect 3010 13572 3066 13628
rect 3066 13572 3070 13628
rect 3006 13568 3070 13572
rect 3086 13628 3150 13632
rect 3086 13572 3090 13628
rect 3090 13572 3146 13628
rect 3146 13572 3150 13628
rect 3086 13568 3150 13572
rect 3166 13628 3230 13632
rect 3166 13572 3170 13628
rect 3170 13572 3226 13628
rect 3226 13572 3230 13628
rect 3166 13568 3230 13572
rect 6874 13628 6938 13632
rect 6874 13572 6878 13628
rect 6878 13572 6934 13628
rect 6934 13572 6938 13628
rect 6874 13568 6938 13572
rect 6954 13628 7018 13632
rect 6954 13572 6958 13628
rect 6958 13572 7014 13628
rect 7014 13572 7018 13628
rect 6954 13568 7018 13572
rect 7034 13628 7098 13632
rect 7034 13572 7038 13628
rect 7038 13572 7094 13628
rect 7094 13572 7098 13628
rect 7034 13568 7098 13572
rect 7114 13628 7178 13632
rect 7114 13572 7118 13628
rect 7118 13572 7174 13628
rect 7174 13572 7178 13628
rect 7114 13568 7178 13572
rect 10822 13628 10886 13632
rect 10822 13572 10826 13628
rect 10826 13572 10882 13628
rect 10882 13572 10886 13628
rect 10822 13568 10886 13572
rect 10902 13628 10966 13632
rect 10902 13572 10906 13628
rect 10906 13572 10962 13628
rect 10962 13572 10966 13628
rect 10902 13568 10966 13572
rect 10982 13628 11046 13632
rect 10982 13572 10986 13628
rect 10986 13572 11042 13628
rect 11042 13572 11046 13628
rect 10982 13568 11046 13572
rect 11062 13628 11126 13632
rect 11062 13572 11066 13628
rect 11066 13572 11122 13628
rect 11122 13572 11126 13628
rect 11062 13568 11126 13572
rect 14770 13628 14834 13632
rect 14770 13572 14774 13628
rect 14774 13572 14830 13628
rect 14830 13572 14834 13628
rect 14770 13568 14834 13572
rect 14850 13628 14914 13632
rect 14850 13572 14854 13628
rect 14854 13572 14910 13628
rect 14910 13572 14914 13628
rect 14850 13568 14914 13572
rect 14930 13628 14994 13632
rect 14930 13572 14934 13628
rect 14934 13572 14990 13628
rect 14990 13572 14994 13628
rect 14930 13568 14994 13572
rect 15010 13628 15074 13632
rect 15010 13572 15014 13628
rect 15014 13572 15070 13628
rect 15070 13572 15074 13628
rect 15010 13568 15074 13572
rect 8708 13364 8772 13428
rect 4900 13084 4964 13088
rect 4900 13028 4904 13084
rect 4904 13028 4960 13084
rect 4960 13028 4964 13084
rect 4900 13024 4964 13028
rect 4980 13084 5044 13088
rect 4980 13028 4984 13084
rect 4984 13028 5040 13084
rect 5040 13028 5044 13084
rect 4980 13024 5044 13028
rect 5060 13084 5124 13088
rect 5060 13028 5064 13084
rect 5064 13028 5120 13084
rect 5120 13028 5124 13084
rect 5060 13024 5124 13028
rect 5140 13084 5204 13088
rect 5140 13028 5144 13084
rect 5144 13028 5200 13084
rect 5200 13028 5204 13084
rect 5140 13024 5204 13028
rect 8848 13084 8912 13088
rect 8848 13028 8852 13084
rect 8852 13028 8908 13084
rect 8908 13028 8912 13084
rect 8848 13024 8912 13028
rect 8928 13084 8992 13088
rect 8928 13028 8932 13084
rect 8932 13028 8988 13084
rect 8988 13028 8992 13084
rect 8928 13024 8992 13028
rect 9008 13084 9072 13088
rect 9008 13028 9012 13084
rect 9012 13028 9068 13084
rect 9068 13028 9072 13084
rect 9008 13024 9072 13028
rect 9088 13084 9152 13088
rect 9088 13028 9092 13084
rect 9092 13028 9148 13084
rect 9148 13028 9152 13084
rect 9088 13024 9152 13028
rect 12796 13084 12860 13088
rect 12796 13028 12800 13084
rect 12800 13028 12856 13084
rect 12856 13028 12860 13084
rect 12796 13024 12860 13028
rect 12876 13084 12940 13088
rect 12876 13028 12880 13084
rect 12880 13028 12936 13084
rect 12936 13028 12940 13084
rect 12876 13024 12940 13028
rect 12956 13084 13020 13088
rect 12956 13028 12960 13084
rect 12960 13028 13016 13084
rect 13016 13028 13020 13084
rect 12956 13024 13020 13028
rect 13036 13084 13100 13088
rect 13036 13028 13040 13084
rect 13040 13028 13096 13084
rect 13096 13028 13100 13084
rect 13036 13024 13100 13028
rect 2926 12540 2990 12544
rect 2926 12484 2930 12540
rect 2930 12484 2986 12540
rect 2986 12484 2990 12540
rect 2926 12480 2990 12484
rect 3006 12540 3070 12544
rect 3006 12484 3010 12540
rect 3010 12484 3066 12540
rect 3066 12484 3070 12540
rect 3006 12480 3070 12484
rect 3086 12540 3150 12544
rect 3086 12484 3090 12540
rect 3090 12484 3146 12540
rect 3146 12484 3150 12540
rect 3086 12480 3150 12484
rect 3166 12540 3230 12544
rect 3166 12484 3170 12540
rect 3170 12484 3226 12540
rect 3226 12484 3230 12540
rect 3166 12480 3230 12484
rect 6874 12540 6938 12544
rect 6874 12484 6878 12540
rect 6878 12484 6934 12540
rect 6934 12484 6938 12540
rect 6874 12480 6938 12484
rect 6954 12540 7018 12544
rect 6954 12484 6958 12540
rect 6958 12484 7014 12540
rect 7014 12484 7018 12540
rect 6954 12480 7018 12484
rect 7034 12540 7098 12544
rect 7034 12484 7038 12540
rect 7038 12484 7094 12540
rect 7094 12484 7098 12540
rect 7034 12480 7098 12484
rect 7114 12540 7178 12544
rect 7114 12484 7118 12540
rect 7118 12484 7174 12540
rect 7174 12484 7178 12540
rect 7114 12480 7178 12484
rect 9260 12412 9324 12476
rect 9444 12472 9508 12476
rect 9444 12416 9494 12472
rect 9494 12416 9508 12472
rect 9444 12412 9508 12416
rect 9812 12276 9876 12340
rect 10822 12540 10886 12544
rect 10822 12484 10826 12540
rect 10826 12484 10882 12540
rect 10882 12484 10886 12540
rect 10822 12480 10886 12484
rect 10902 12540 10966 12544
rect 10902 12484 10906 12540
rect 10906 12484 10962 12540
rect 10962 12484 10966 12540
rect 10902 12480 10966 12484
rect 10982 12540 11046 12544
rect 10982 12484 10986 12540
rect 10986 12484 11042 12540
rect 11042 12484 11046 12540
rect 10982 12480 11046 12484
rect 11062 12540 11126 12544
rect 11062 12484 11066 12540
rect 11066 12484 11122 12540
rect 11122 12484 11126 12540
rect 11062 12480 11126 12484
rect 14770 12540 14834 12544
rect 14770 12484 14774 12540
rect 14774 12484 14830 12540
rect 14830 12484 14834 12540
rect 14770 12480 14834 12484
rect 14850 12540 14914 12544
rect 14850 12484 14854 12540
rect 14854 12484 14910 12540
rect 14910 12484 14914 12540
rect 14850 12480 14914 12484
rect 14930 12540 14994 12544
rect 14930 12484 14934 12540
rect 14934 12484 14990 12540
rect 14990 12484 14994 12540
rect 14930 12480 14994 12484
rect 15010 12540 15074 12544
rect 15010 12484 15014 12540
rect 15014 12484 15070 12540
rect 15070 12484 15074 12540
rect 15010 12480 15074 12484
rect 8524 12064 8588 12068
rect 8524 12008 8574 12064
rect 8574 12008 8588 12064
rect 8524 12004 8588 12008
rect 9260 12004 9324 12068
rect 4900 11996 4964 12000
rect 4900 11940 4904 11996
rect 4904 11940 4960 11996
rect 4960 11940 4964 11996
rect 4900 11936 4964 11940
rect 4980 11996 5044 12000
rect 4980 11940 4984 11996
rect 4984 11940 5040 11996
rect 5040 11940 5044 11996
rect 4980 11936 5044 11940
rect 5060 11996 5124 12000
rect 5060 11940 5064 11996
rect 5064 11940 5120 11996
rect 5120 11940 5124 11996
rect 5060 11936 5124 11940
rect 5140 11996 5204 12000
rect 5140 11940 5144 11996
rect 5144 11940 5200 11996
rect 5200 11940 5204 11996
rect 5140 11936 5204 11940
rect 8848 11996 8912 12000
rect 8848 11940 8852 11996
rect 8852 11940 8908 11996
rect 8908 11940 8912 11996
rect 8848 11936 8912 11940
rect 8928 11996 8992 12000
rect 8928 11940 8932 11996
rect 8932 11940 8988 11996
rect 8988 11940 8992 11996
rect 8928 11936 8992 11940
rect 9008 11996 9072 12000
rect 9008 11940 9012 11996
rect 9012 11940 9068 11996
rect 9068 11940 9072 11996
rect 9008 11936 9072 11940
rect 9088 11996 9152 12000
rect 9088 11940 9092 11996
rect 9092 11940 9148 11996
rect 9148 11940 9152 11996
rect 9088 11936 9152 11940
rect 12796 11996 12860 12000
rect 12796 11940 12800 11996
rect 12800 11940 12856 11996
rect 12856 11940 12860 11996
rect 12796 11936 12860 11940
rect 12876 11996 12940 12000
rect 12876 11940 12880 11996
rect 12880 11940 12936 11996
rect 12936 11940 12940 11996
rect 12876 11936 12940 11940
rect 12956 11996 13020 12000
rect 12956 11940 12960 11996
rect 12960 11940 13016 11996
rect 13016 11940 13020 11996
rect 12956 11936 13020 11940
rect 13036 11996 13100 12000
rect 13036 11940 13040 11996
rect 13040 11940 13096 11996
rect 13096 11940 13100 11996
rect 13036 11936 13100 11940
rect 3556 11732 3620 11796
rect 8708 11732 8772 11796
rect 10548 11732 10612 11796
rect 3740 11460 3804 11524
rect 2926 11452 2990 11456
rect 2926 11396 2930 11452
rect 2930 11396 2986 11452
rect 2986 11396 2990 11452
rect 2926 11392 2990 11396
rect 3006 11452 3070 11456
rect 3006 11396 3010 11452
rect 3010 11396 3066 11452
rect 3066 11396 3070 11452
rect 3006 11392 3070 11396
rect 3086 11452 3150 11456
rect 3086 11396 3090 11452
rect 3090 11396 3146 11452
rect 3146 11396 3150 11452
rect 3086 11392 3150 11396
rect 3166 11452 3230 11456
rect 3166 11396 3170 11452
rect 3170 11396 3226 11452
rect 3226 11396 3230 11452
rect 3166 11392 3230 11396
rect 6874 11452 6938 11456
rect 6874 11396 6878 11452
rect 6878 11396 6934 11452
rect 6934 11396 6938 11452
rect 6874 11392 6938 11396
rect 6954 11452 7018 11456
rect 6954 11396 6958 11452
rect 6958 11396 7014 11452
rect 7014 11396 7018 11452
rect 6954 11392 7018 11396
rect 7034 11452 7098 11456
rect 7034 11396 7038 11452
rect 7038 11396 7094 11452
rect 7094 11396 7098 11452
rect 7034 11392 7098 11396
rect 7114 11452 7178 11456
rect 7114 11396 7118 11452
rect 7118 11396 7174 11452
rect 7174 11396 7178 11452
rect 7114 11392 7178 11396
rect 10822 11452 10886 11456
rect 10822 11396 10826 11452
rect 10826 11396 10882 11452
rect 10882 11396 10886 11452
rect 10822 11392 10886 11396
rect 10902 11452 10966 11456
rect 10902 11396 10906 11452
rect 10906 11396 10962 11452
rect 10962 11396 10966 11452
rect 10902 11392 10966 11396
rect 10982 11452 11046 11456
rect 10982 11396 10986 11452
rect 10986 11396 11042 11452
rect 11042 11396 11046 11452
rect 10982 11392 11046 11396
rect 11062 11452 11126 11456
rect 11062 11396 11066 11452
rect 11066 11396 11122 11452
rect 11122 11396 11126 11452
rect 11062 11392 11126 11396
rect 14770 11452 14834 11456
rect 14770 11396 14774 11452
rect 14774 11396 14830 11452
rect 14830 11396 14834 11452
rect 14770 11392 14834 11396
rect 14850 11452 14914 11456
rect 14850 11396 14854 11452
rect 14854 11396 14910 11452
rect 14910 11396 14914 11452
rect 14850 11392 14914 11396
rect 14930 11452 14994 11456
rect 14930 11396 14934 11452
rect 14934 11396 14990 11452
rect 14990 11396 14994 11452
rect 14930 11392 14994 11396
rect 15010 11452 15074 11456
rect 15010 11396 15014 11452
rect 15014 11396 15070 11452
rect 15070 11396 15074 11452
rect 15010 11392 15074 11396
rect 2636 11052 2700 11116
rect 5948 11052 6012 11116
rect 4900 10908 4964 10912
rect 4900 10852 4904 10908
rect 4904 10852 4960 10908
rect 4960 10852 4964 10908
rect 4900 10848 4964 10852
rect 4980 10908 5044 10912
rect 4980 10852 4984 10908
rect 4984 10852 5040 10908
rect 5040 10852 5044 10908
rect 4980 10848 5044 10852
rect 5060 10908 5124 10912
rect 5060 10852 5064 10908
rect 5064 10852 5120 10908
rect 5120 10852 5124 10908
rect 5060 10848 5124 10852
rect 5140 10908 5204 10912
rect 5140 10852 5144 10908
rect 5144 10852 5200 10908
rect 5200 10852 5204 10908
rect 5140 10848 5204 10852
rect 8848 10908 8912 10912
rect 8848 10852 8852 10908
rect 8852 10852 8908 10908
rect 8908 10852 8912 10908
rect 8848 10848 8912 10852
rect 8928 10908 8992 10912
rect 8928 10852 8932 10908
rect 8932 10852 8988 10908
rect 8988 10852 8992 10908
rect 8928 10848 8992 10852
rect 9008 10908 9072 10912
rect 9008 10852 9012 10908
rect 9012 10852 9068 10908
rect 9068 10852 9072 10908
rect 9008 10848 9072 10852
rect 9088 10908 9152 10912
rect 9088 10852 9092 10908
rect 9092 10852 9148 10908
rect 9148 10852 9152 10908
rect 9088 10848 9152 10852
rect 12796 10908 12860 10912
rect 12796 10852 12800 10908
rect 12800 10852 12856 10908
rect 12856 10852 12860 10908
rect 12796 10848 12860 10852
rect 12876 10908 12940 10912
rect 12876 10852 12880 10908
rect 12880 10852 12936 10908
rect 12936 10852 12940 10908
rect 12876 10848 12940 10852
rect 12956 10908 13020 10912
rect 12956 10852 12960 10908
rect 12960 10852 13016 10908
rect 13016 10852 13020 10908
rect 12956 10848 13020 10852
rect 13036 10908 13100 10912
rect 13036 10852 13040 10908
rect 13040 10852 13096 10908
rect 13096 10852 13100 10908
rect 13036 10848 13100 10852
rect 9812 10780 9876 10844
rect 8156 10644 8220 10708
rect 7972 10372 8036 10436
rect 2926 10364 2990 10368
rect 2926 10308 2930 10364
rect 2930 10308 2986 10364
rect 2986 10308 2990 10364
rect 2926 10304 2990 10308
rect 3006 10364 3070 10368
rect 3006 10308 3010 10364
rect 3010 10308 3066 10364
rect 3066 10308 3070 10364
rect 3006 10304 3070 10308
rect 3086 10364 3150 10368
rect 3086 10308 3090 10364
rect 3090 10308 3146 10364
rect 3146 10308 3150 10364
rect 3086 10304 3150 10308
rect 3166 10364 3230 10368
rect 3166 10308 3170 10364
rect 3170 10308 3226 10364
rect 3226 10308 3230 10364
rect 3166 10304 3230 10308
rect 6874 10364 6938 10368
rect 6874 10308 6878 10364
rect 6878 10308 6934 10364
rect 6934 10308 6938 10364
rect 6874 10304 6938 10308
rect 6954 10364 7018 10368
rect 6954 10308 6958 10364
rect 6958 10308 7014 10364
rect 7014 10308 7018 10364
rect 6954 10304 7018 10308
rect 7034 10364 7098 10368
rect 7034 10308 7038 10364
rect 7038 10308 7094 10364
rect 7094 10308 7098 10364
rect 7034 10304 7098 10308
rect 7114 10364 7178 10368
rect 7114 10308 7118 10364
rect 7118 10308 7174 10364
rect 7174 10308 7178 10364
rect 7114 10304 7178 10308
rect 7420 10236 7484 10300
rect 10822 10364 10886 10368
rect 10822 10308 10826 10364
rect 10826 10308 10882 10364
rect 10882 10308 10886 10364
rect 10822 10304 10886 10308
rect 10902 10364 10966 10368
rect 10902 10308 10906 10364
rect 10906 10308 10962 10364
rect 10962 10308 10966 10364
rect 10902 10304 10966 10308
rect 10982 10364 11046 10368
rect 10982 10308 10986 10364
rect 10986 10308 11042 10364
rect 11042 10308 11046 10364
rect 10982 10304 11046 10308
rect 11062 10364 11126 10368
rect 11062 10308 11066 10364
rect 11066 10308 11122 10364
rect 11122 10308 11126 10364
rect 11062 10304 11126 10308
rect 14770 10364 14834 10368
rect 14770 10308 14774 10364
rect 14774 10308 14830 10364
rect 14830 10308 14834 10364
rect 14770 10304 14834 10308
rect 14850 10364 14914 10368
rect 14850 10308 14854 10364
rect 14854 10308 14910 10364
rect 14910 10308 14914 10364
rect 14850 10304 14914 10308
rect 14930 10364 14994 10368
rect 14930 10308 14934 10364
rect 14934 10308 14990 10364
rect 14990 10308 14994 10364
rect 14930 10304 14994 10308
rect 15010 10364 15074 10368
rect 15010 10308 15014 10364
rect 15014 10308 15070 10364
rect 15070 10308 15074 10364
rect 15010 10304 15074 10308
rect 2636 9964 2700 10028
rect 4900 9820 4964 9824
rect 4900 9764 4904 9820
rect 4904 9764 4960 9820
rect 4960 9764 4964 9820
rect 4900 9760 4964 9764
rect 4980 9820 5044 9824
rect 4980 9764 4984 9820
rect 4984 9764 5040 9820
rect 5040 9764 5044 9820
rect 4980 9760 5044 9764
rect 5060 9820 5124 9824
rect 5060 9764 5064 9820
rect 5064 9764 5120 9820
rect 5120 9764 5124 9820
rect 5060 9760 5124 9764
rect 5140 9820 5204 9824
rect 5140 9764 5144 9820
rect 5144 9764 5200 9820
rect 5200 9764 5204 9820
rect 5140 9760 5204 9764
rect 8848 9820 8912 9824
rect 8848 9764 8852 9820
rect 8852 9764 8908 9820
rect 8908 9764 8912 9820
rect 8848 9760 8912 9764
rect 8928 9820 8992 9824
rect 8928 9764 8932 9820
rect 8932 9764 8988 9820
rect 8988 9764 8992 9820
rect 8928 9760 8992 9764
rect 9008 9820 9072 9824
rect 9008 9764 9012 9820
rect 9012 9764 9068 9820
rect 9068 9764 9072 9820
rect 9008 9760 9072 9764
rect 9088 9820 9152 9824
rect 9088 9764 9092 9820
rect 9092 9764 9148 9820
rect 9148 9764 9152 9820
rect 9088 9760 9152 9764
rect 12796 9820 12860 9824
rect 12796 9764 12800 9820
rect 12800 9764 12856 9820
rect 12856 9764 12860 9820
rect 12796 9760 12860 9764
rect 12876 9820 12940 9824
rect 12876 9764 12880 9820
rect 12880 9764 12936 9820
rect 12936 9764 12940 9820
rect 12876 9760 12940 9764
rect 12956 9820 13020 9824
rect 12956 9764 12960 9820
rect 12960 9764 13016 9820
rect 13016 9764 13020 9820
rect 12956 9760 13020 9764
rect 13036 9820 13100 9824
rect 13036 9764 13040 9820
rect 13040 9764 13096 9820
rect 13096 9764 13100 9820
rect 13036 9760 13100 9764
rect 9628 9692 9692 9756
rect 4660 9556 4724 9620
rect 9996 9480 10060 9484
rect 9996 9424 10010 9480
rect 10010 9424 10060 9480
rect 9996 9420 10060 9424
rect 2926 9276 2990 9280
rect 2926 9220 2930 9276
rect 2930 9220 2986 9276
rect 2986 9220 2990 9276
rect 2926 9216 2990 9220
rect 3006 9276 3070 9280
rect 3006 9220 3010 9276
rect 3010 9220 3066 9276
rect 3066 9220 3070 9276
rect 3006 9216 3070 9220
rect 3086 9276 3150 9280
rect 3086 9220 3090 9276
rect 3090 9220 3146 9276
rect 3146 9220 3150 9276
rect 3086 9216 3150 9220
rect 3166 9276 3230 9280
rect 3166 9220 3170 9276
rect 3170 9220 3226 9276
rect 3226 9220 3230 9276
rect 3166 9216 3230 9220
rect 6874 9276 6938 9280
rect 6874 9220 6878 9276
rect 6878 9220 6934 9276
rect 6934 9220 6938 9276
rect 6874 9216 6938 9220
rect 6954 9276 7018 9280
rect 6954 9220 6958 9276
rect 6958 9220 7014 9276
rect 7014 9220 7018 9276
rect 6954 9216 7018 9220
rect 7034 9276 7098 9280
rect 7034 9220 7038 9276
rect 7038 9220 7094 9276
rect 7094 9220 7098 9276
rect 7034 9216 7098 9220
rect 7114 9276 7178 9280
rect 7114 9220 7118 9276
rect 7118 9220 7174 9276
rect 7174 9220 7178 9276
rect 7114 9216 7178 9220
rect 10822 9276 10886 9280
rect 10822 9220 10826 9276
rect 10826 9220 10882 9276
rect 10882 9220 10886 9276
rect 10822 9216 10886 9220
rect 10902 9276 10966 9280
rect 10902 9220 10906 9276
rect 10906 9220 10962 9276
rect 10962 9220 10966 9276
rect 10902 9216 10966 9220
rect 10982 9276 11046 9280
rect 10982 9220 10986 9276
rect 10986 9220 11042 9276
rect 11042 9220 11046 9276
rect 10982 9216 11046 9220
rect 11062 9276 11126 9280
rect 11062 9220 11066 9276
rect 11066 9220 11122 9276
rect 11122 9220 11126 9276
rect 11062 9216 11126 9220
rect 14770 9276 14834 9280
rect 14770 9220 14774 9276
rect 14774 9220 14830 9276
rect 14830 9220 14834 9276
rect 14770 9216 14834 9220
rect 14850 9276 14914 9280
rect 14850 9220 14854 9276
rect 14854 9220 14910 9276
rect 14910 9220 14914 9276
rect 14850 9216 14914 9220
rect 14930 9276 14994 9280
rect 14930 9220 14934 9276
rect 14934 9220 14990 9276
rect 14990 9220 14994 9276
rect 14930 9216 14994 9220
rect 15010 9276 15074 9280
rect 15010 9220 15014 9276
rect 15014 9220 15070 9276
rect 15070 9220 15074 9276
rect 15010 9216 15074 9220
rect 9260 9148 9324 9212
rect 10180 9148 10244 9212
rect 10364 9148 10428 9212
rect 8340 8876 8404 8940
rect 6684 8740 6748 8804
rect 9444 8740 9508 8804
rect 4900 8732 4964 8736
rect 4900 8676 4904 8732
rect 4904 8676 4960 8732
rect 4960 8676 4964 8732
rect 4900 8672 4964 8676
rect 4980 8732 5044 8736
rect 4980 8676 4984 8732
rect 4984 8676 5040 8732
rect 5040 8676 5044 8732
rect 4980 8672 5044 8676
rect 5060 8732 5124 8736
rect 5060 8676 5064 8732
rect 5064 8676 5120 8732
rect 5120 8676 5124 8732
rect 5060 8672 5124 8676
rect 5140 8732 5204 8736
rect 5140 8676 5144 8732
rect 5144 8676 5200 8732
rect 5200 8676 5204 8732
rect 5140 8672 5204 8676
rect 8848 8732 8912 8736
rect 8848 8676 8852 8732
rect 8852 8676 8908 8732
rect 8908 8676 8912 8732
rect 8848 8672 8912 8676
rect 8928 8732 8992 8736
rect 8928 8676 8932 8732
rect 8932 8676 8988 8732
rect 8988 8676 8992 8732
rect 8928 8672 8992 8676
rect 9008 8732 9072 8736
rect 9008 8676 9012 8732
rect 9012 8676 9068 8732
rect 9068 8676 9072 8732
rect 9008 8672 9072 8676
rect 9088 8732 9152 8736
rect 9088 8676 9092 8732
rect 9092 8676 9148 8732
rect 9148 8676 9152 8732
rect 9088 8672 9152 8676
rect 12796 8732 12860 8736
rect 12796 8676 12800 8732
rect 12800 8676 12856 8732
rect 12856 8676 12860 8732
rect 12796 8672 12860 8676
rect 12876 8732 12940 8736
rect 12876 8676 12880 8732
rect 12880 8676 12936 8732
rect 12936 8676 12940 8732
rect 12876 8672 12940 8676
rect 12956 8732 13020 8736
rect 12956 8676 12960 8732
rect 12960 8676 13016 8732
rect 13016 8676 13020 8732
rect 12956 8672 13020 8676
rect 13036 8732 13100 8736
rect 13036 8676 13040 8732
rect 13040 8676 13096 8732
rect 13096 8676 13100 8732
rect 13036 8672 13100 8676
rect 9260 8604 9324 8668
rect 5580 8332 5644 8396
rect 7420 8332 7484 8396
rect 8708 8332 8772 8396
rect 9444 8332 9508 8396
rect 9812 8332 9876 8396
rect 11284 8392 11348 8396
rect 11284 8336 11298 8392
rect 11298 8336 11348 8392
rect 11284 8332 11348 8336
rect 2926 8188 2990 8192
rect 2926 8132 2930 8188
rect 2930 8132 2986 8188
rect 2986 8132 2990 8188
rect 2926 8128 2990 8132
rect 3006 8188 3070 8192
rect 3006 8132 3010 8188
rect 3010 8132 3066 8188
rect 3066 8132 3070 8188
rect 3006 8128 3070 8132
rect 3086 8188 3150 8192
rect 3086 8132 3090 8188
rect 3090 8132 3146 8188
rect 3146 8132 3150 8188
rect 3086 8128 3150 8132
rect 3166 8188 3230 8192
rect 3166 8132 3170 8188
rect 3170 8132 3226 8188
rect 3226 8132 3230 8188
rect 3166 8128 3230 8132
rect 6874 8188 6938 8192
rect 6874 8132 6878 8188
rect 6878 8132 6934 8188
rect 6934 8132 6938 8188
rect 6874 8128 6938 8132
rect 6954 8188 7018 8192
rect 6954 8132 6958 8188
rect 6958 8132 7014 8188
rect 7014 8132 7018 8188
rect 6954 8128 7018 8132
rect 7034 8188 7098 8192
rect 7034 8132 7038 8188
rect 7038 8132 7094 8188
rect 7094 8132 7098 8188
rect 7034 8128 7098 8132
rect 7114 8188 7178 8192
rect 7114 8132 7118 8188
rect 7118 8132 7174 8188
rect 7174 8132 7178 8188
rect 7114 8128 7178 8132
rect 10822 8188 10886 8192
rect 10822 8132 10826 8188
rect 10826 8132 10882 8188
rect 10882 8132 10886 8188
rect 10822 8128 10886 8132
rect 10902 8188 10966 8192
rect 10902 8132 10906 8188
rect 10906 8132 10962 8188
rect 10962 8132 10966 8188
rect 10902 8128 10966 8132
rect 10982 8188 11046 8192
rect 10982 8132 10986 8188
rect 10986 8132 11042 8188
rect 11042 8132 11046 8188
rect 10982 8128 11046 8132
rect 11062 8188 11126 8192
rect 11062 8132 11066 8188
rect 11066 8132 11122 8188
rect 11122 8132 11126 8188
rect 11062 8128 11126 8132
rect 14770 8188 14834 8192
rect 14770 8132 14774 8188
rect 14774 8132 14830 8188
rect 14830 8132 14834 8188
rect 14770 8128 14834 8132
rect 14850 8188 14914 8192
rect 14850 8132 14854 8188
rect 14854 8132 14910 8188
rect 14910 8132 14914 8188
rect 14850 8128 14914 8132
rect 14930 8188 14994 8192
rect 14930 8132 14934 8188
rect 14934 8132 14990 8188
rect 14990 8132 14994 8188
rect 14930 8128 14994 8132
rect 15010 8188 15074 8192
rect 15010 8132 15014 8188
rect 15014 8132 15070 8188
rect 15070 8132 15074 8188
rect 15010 8128 15074 8132
rect 5764 8120 5828 8124
rect 5764 8064 5778 8120
rect 5778 8064 5828 8120
rect 5764 8060 5828 8064
rect 6132 8120 6196 8124
rect 6132 8064 6182 8120
rect 6182 8064 6196 8120
rect 6132 8060 6196 8064
rect 6316 8120 6380 8124
rect 6316 8064 6366 8120
rect 6366 8064 6380 8120
rect 6316 8060 6380 8064
rect 10548 8060 10612 8124
rect 10364 7788 10428 7852
rect 4900 7644 4964 7648
rect 4900 7588 4904 7644
rect 4904 7588 4960 7644
rect 4960 7588 4964 7644
rect 4900 7584 4964 7588
rect 4980 7644 5044 7648
rect 4980 7588 4984 7644
rect 4984 7588 5040 7644
rect 5040 7588 5044 7644
rect 4980 7584 5044 7588
rect 5060 7644 5124 7648
rect 5060 7588 5064 7644
rect 5064 7588 5120 7644
rect 5120 7588 5124 7644
rect 5060 7584 5124 7588
rect 5140 7644 5204 7648
rect 5140 7588 5144 7644
rect 5144 7588 5200 7644
rect 5200 7588 5204 7644
rect 5140 7584 5204 7588
rect 10180 7652 10244 7716
rect 8848 7644 8912 7648
rect 8848 7588 8852 7644
rect 8852 7588 8908 7644
rect 8908 7588 8912 7644
rect 8848 7584 8912 7588
rect 8928 7644 8992 7648
rect 8928 7588 8932 7644
rect 8932 7588 8988 7644
rect 8988 7588 8992 7644
rect 8928 7584 8992 7588
rect 9008 7644 9072 7648
rect 9008 7588 9012 7644
rect 9012 7588 9068 7644
rect 9068 7588 9072 7644
rect 9008 7584 9072 7588
rect 9088 7644 9152 7648
rect 9088 7588 9092 7644
rect 9092 7588 9148 7644
rect 9148 7588 9152 7644
rect 9088 7584 9152 7588
rect 12796 7644 12860 7648
rect 12796 7588 12800 7644
rect 12800 7588 12856 7644
rect 12856 7588 12860 7644
rect 12796 7584 12860 7588
rect 12876 7644 12940 7648
rect 12876 7588 12880 7644
rect 12880 7588 12936 7644
rect 12936 7588 12940 7644
rect 12876 7584 12940 7588
rect 12956 7644 13020 7648
rect 12956 7588 12960 7644
rect 12960 7588 13016 7644
rect 13016 7588 13020 7644
rect 12956 7584 13020 7588
rect 13036 7644 13100 7648
rect 13036 7588 13040 7644
rect 13040 7588 13096 7644
rect 13096 7588 13100 7644
rect 13036 7584 13100 7588
rect 5948 7576 6012 7580
rect 5948 7520 5962 7576
rect 5962 7520 6012 7576
rect 5948 7516 6012 7520
rect 9996 7516 10060 7580
rect 6132 7108 6196 7172
rect 6500 7108 6564 7172
rect 2926 7100 2990 7104
rect 2926 7044 2930 7100
rect 2930 7044 2986 7100
rect 2986 7044 2990 7100
rect 2926 7040 2990 7044
rect 3006 7100 3070 7104
rect 3006 7044 3010 7100
rect 3010 7044 3066 7100
rect 3066 7044 3070 7100
rect 3006 7040 3070 7044
rect 3086 7100 3150 7104
rect 3086 7044 3090 7100
rect 3090 7044 3146 7100
rect 3146 7044 3150 7100
rect 3086 7040 3150 7044
rect 3166 7100 3230 7104
rect 3166 7044 3170 7100
rect 3170 7044 3226 7100
rect 3226 7044 3230 7100
rect 3166 7040 3230 7044
rect 6874 7100 6938 7104
rect 6874 7044 6878 7100
rect 6878 7044 6934 7100
rect 6934 7044 6938 7100
rect 6874 7040 6938 7044
rect 6954 7100 7018 7104
rect 6954 7044 6958 7100
rect 6958 7044 7014 7100
rect 7014 7044 7018 7100
rect 6954 7040 7018 7044
rect 7034 7100 7098 7104
rect 7034 7044 7038 7100
rect 7038 7044 7094 7100
rect 7094 7044 7098 7100
rect 7034 7040 7098 7044
rect 7114 7100 7178 7104
rect 7114 7044 7118 7100
rect 7118 7044 7174 7100
rect 7174 7044 7178 7100
rect 7114 7040 7178 7044
rect 4108 7032 4172 7036
rect 4108 6976 4158 7032
rect 4158 6976 4172 7032
rect 4108 6972 4172 6976
rect 10822 7100 10886 7104
rect 10822 7044 10826 7100
rect 10826 7044 10882 7100
rect 10882 7044 10886 7100
rect 10822 7040 10886 7044
rect 10902 7100 10966 7104
rect 10902 7044 10906 7100
rect 10906 7044 10962 7100
rect 10962 7044 10966 7100
rect 10902 7040 10966 7044
rect 10982 7100 11046 7104
rect 10982 7044 10986 7100
rect 10986 7044 11042 7100
rect 11042 7044 11046 7100
rect 10982 7040 11046 7044
rect 11062 7100 11126 7104
rect 11062 7044 11066 7100
rect 11066 7044 11122 7100
rect 11122 7044 11126 7100
rect 11062 7040 11126 7044
rect 14770 7100 14834 7104
rect 14770 7044 14774 7100
rect 14774 7044 14830 7100
rect 14830 7044 14834 7100
rect 14770 7040 14834 7044
rect 14850 7100 14914 7104
rect 14850 7044 14854 7100
rect 14854 7044 14910 7100
rect 14910 7044 14914 7100
rect 14850 7040 14914 7044
rect 14930 7100 14994 7104
rect 14930 7044 14934 7100
rect 14934 7044 14990 7100
rect 14990 7044 14994 7100
rect 14930 7040 14994 7044
rect 15010 7100 15074 7104
rect 15010 7044 15014 7100
rect 15014 7044 15070 7100
rect 15070 7044 15074 7100
rect 15010 7040 15074 7044
rect 6316 6896 6380 6900
rect 6316 6840 6366 6896
rect 6366 6840 6380 6896
rect 6316 6836 6380 6840
rect 5764 6624 5828 6628
rect 5764 6568 5814 6624
rect 5814 6568 5828 6624
rect 5764 6564 5828 6568
rect 8156 6564 8220 6628
rect 4900 6556 4964 6560
rect 4900 6500 4904 6556
rect 4904 6500 4960 6556
rect 4960 6500 4964 6556
rect 4900 6496 4964 6500
rect 4980 6556 5044 6560
rect 4980 6500 4984 6556
rect 4984 6500 5040 6556
rect 5040 6500 5044 6556
rect 4980 6496 5044 6500
rect 5060 6556 5124 6560
rect 5060 6500 5064 6556
rect 5064 6500 5120 6556
rect 5120 6500 5124 6556
rect 5060 6496 5124 6500
rect 5140 6556 5204 6560
rect 5140 6500 5144 6556
rect 5144 6500 5200 6556
rect 5200 6500 5204 6556
rect 5140 6496 5204 6500
rect 8848 6556 8912 6560
rect 8848 6500 8852 6556
rect 8852 6500 8908 6556
rect 8908 6500 8912 6556
rect 8848 6496 8912 6500
rect 8928 6556 8992 6560
rect 8928 6500 8932 6556
rect 8932 6500 8988 6556
rect 8988 6500 8992 6556
rect 8928 6496 8992 6500
rect 9008 6556 9072 6560
rect 9008 6500 9012 6556
rect 9012 6500 9068 6556
rect 9068 6500 9072 6556
rect 9008 6496 9072 6500
rect 9088 6556 9152 6560
rect 9088 6500 9092 6556
rect 9092 6500 9148 6556
rect 9148 6500 9152 6556
rect 9088 6496 9152 6500
rect 12796 6556 12860 6560
rect 12796 6500 12800 6556
rect 12800 6500 12856 6556
rect 12856 6500 12860 6556
rect 12796 6496 12860 6500
rect 12876 6556 12940 6560
rect 12876 6500 12880 6556
rect 12880 6500 12936 6556
rect 12936 6500 12940 6556
rect 12876 6496 12940 6500
rect 12956 6556 13020 6560
rect 12956 6500 12960 6556
rect 12960 6500 13016 6556
rect 13016 6500 13020 6556
rect 12956 6496 13020 6500
rect 13036 6556 13100 6560
rect 13036 6500 13040 6556
rect 13040 6500 13096 6556
rect 13096 6500 13100 6556
rect 13036 6496 13100 6500
rect 6684 6428 6748 6492
rect 7972 6428 8036 6492
rect 2926 6012 2990 6016
rect 2926 5956 2930 6012
rect 2930 5956 2986 6012
rect 2986 5956 2990 6012
rect 2926 5952 2990 5956
rect 3006 6012 3070 6016
rect 3006 5956 3010 6012
rect 3010 5956 3066 6012
rect 3066 5956 3070 6012
rect 3006 5952 3070 5956
rect 3086 6012 3150 6016
rect 3086 5956 3090 6012
rect 3090 5956 3146 6012
rect 3146 5956 3150 6012
rect 3086 5952 3150 5956
rect 3166 6012 3230 6016
rect 3166 5956 3170 6012
rect 3170 5956 3226 6012
rect 3226 5956 3230 6012
rect 3166 5952 3230 5956
rect 6874 6012 6938 6016
rect 6874 5956 6878 6012
rect 6878 5956 6934 6012
rect 6934 5956 6938 6012
rect 6874 5952 6938 5956
rect 6954 6012 7018 6016
rect 6954 5956 6958 6012
rect 6958 5956 7014 6012
rect 7014 5956 7018 6012
rect 6954 5952 7018 5956
rect 7034 6012 7098 6016
rect 7034 5956 7038 6012
rect 7038 5956 7094 6012
rect 7094 5956 7098 6012
rect 7034 5952 7098 5956
rect 7114 6012 7178 6016
rect 7114 5956 7118 6012
rect 7118 5956 7174 6012
rect 7174 5956 7178 6012
rect 7114 5952 7178 5956
rect 10822 6012 10886 6016
rect 10822 5956 10826 6012
rect 10826 5956 10882 6012
rect 10882 5956 10886 6012
rect 10822 5952 10886 5956
rect 10902 6012 10966 6016
rect 10902 5956 10906 6012
rect 10906 5956 10962 6012
rect 10962 5956 10966 6012
rect 10902 5952 10966 5956
rect 10982 6012 11046 6016
rect 10982 5956 10986 6012
rect 10986 5956 11042 6012
rect 11042 5956 11046 6012
rect 10982 5952 11046 5956
rect 11062 6012 11126 6016
rect 11062 5956 11066 6012
rect 11066 5956 11122 6012
rect 11122 5956 11126 6012
rect 11062 5952 11126 5956
rect 14770 6012 14834 6016
rect 14770 5956 14774 6012
rect 14774 5956 14830 6012
rect 14830 5956 14834 6012
rect 14770 5952 14834 5956
rect 14850 6012 14914 6016
rect 14850 5956 14854 6012
rect 14854 5956 14910 6012
rect 14910 5956 14914 6012
rect 14850 5952 14914 5956
rect 14930 6012 14994 6016
rect 14930 5956 14934 6012
rect 14934 5956 14990 6012
rect 14990 5956 14994 6012
rect 14930 5952 14994 5956
rect 15010 6012 15074 6016
rect 15010 5956 15014 6012
rect 15014 5956 15070 6012
rect 15070 5956 15074 6012
rect 15010 5952 15074 5956
rect 9628 5748 9692 5812
rect 4900 5468 4964 5472
rect 4900 5412 4904 5468
rect 4904 5412 4960 5468
rect 4960 5412 4964 5468
rect 4900 5408 4964 5412
rect 4980 5468 5044 5472
rect 4980 5412 4984 5468
rect 4984 5412 5040 5468
rect 5040 5412 5044 5468
rect 4980 5408 5044 5412
rect 5060 5468 5124 5472
rect 5060 5412 5064 5468
rect 5064 5412 5120 5468
rect 5120 5412 5124 5468
rect 5060 5408 5124 5412
rect 5140 5468 5204 5472
rect 5140 5412 5144 5468
rect 5144 5412 5200 5468
rect 5200 5412 5204 5468
rect 5140 5408 5204 5412
rect 8848 5468 8912 5472
rect 8848 5412 8852 5468
rect 8852 5412 8908 5468
rect 8908 5412 8912 5468
rect 8848 5408 8912 5412
rect 8928 5468 8992 5472
rect 8928 5412 8932 5468
rect 8932 5412 8988 5468
rect 8988 5412 8992 5468
rect 8928 5408 8992 5412
rect 9008 5468 9072 5472
rect 9008 5412 9012 5468
rect 9012 5412 9068 5468
rect 9068 5412 9072 5468
rect 9008 5408 9072 5412
rect 9088 5468 9152 5472
rect 9088 5412 9092 5468
rect 9092 5412 9148 5468
rect 9148 5412 9152 5468
rect 9088 5408 9152 5412
rect 12796 5468 12860 5472
rect 12796 5412 12800 5468
rect 12800 5412 12856 5468
rect 12856 5412 12860 5468
rect 12796 5408 12860 5412
rect 12876 5468 12940 5472
rect 12876 5412 12880 5468
rect 12880 5412 12936 5468
rect 12936 5412 12940 5468
rect 12876 5408 12940 5412
rect 12956 5468 13020 5472
rect 12956 5412 12960 5468
rect 12960 5412 13016 5468
rect 13016 5412 13020 5468
rect 12956 5408 13020 5412
rect 13036 5468 13100 5472
rect 13036 5412 13040 5468
rect 13040 5412 13096 5468
rect 13096 5412 13100 5468
rect 13036 5408 13100 5412
rect 3556 5340 3620 5404
rect 5396 5400 5460 5404
rect 5396 5344 5410 5400
rect 5410 5344 5460 5400
rect 5396 5340 5460 5344
rect 8524 5400 8588 5404
rect 8524 5344 8538 5400
rect 8538 5344 8588 5400
rect 8524 5340 8588 5344
rect 7420 5204 7484 5268
rect 11284 5068 11348 5132
rect 4660 4992 4724 4996
rect 4660 4936 4710 4992
rect 4710 4936 4724 4992
rect 4660 4932 4724 4936
rect 2926 4924 2990 4928
rect 2926 4868 2930 4924
rect 2930 4868 2986 4924
rect 2986 4868 2990 4924
rect 2926 4864 2990 4868
rect 3006 4924 3070 4928
rect 3006 4868 3010 4924
rect 3010 4868 3066 4924
rect 3066 4868 3070 4924
rect 3006 4864 3070 4868
rect 3086 4924 3150 4928
rect 3086 4868 3090 4924
rect 3090 4868 3146 4924
rect 3146 4868 3150 4924
rect 3086 4864 3150 4868
rect 3166 4924 3230 4928
rect 3166 4868 3170 4924
rect 3170 4868 3226 4924
rect 3226 4868 3230 4924
rect 3166 4864 3230 4868
rect 6874 4924 6938 4928
rect 6874 4868 6878 4924
rect 6878 4868 6934 4924
rect 6934 4868 6938 4924
rect 6874 4864 6938 4868
rect 6954 4924 7018 4928
rect 6954 4868 6958 4924
rect 6958 4868 7014 4924
rect 7014 4868 7018 4924
rect 6954 4864 7018 4868
rect 7034 4924 7098 4928
rect 7034 4868 7038 4924
rect 7038 4868 7094 4924
rect 7094 4868 7098 4924
rect 7034 4864 7098 4868
rect 7114 4924 7178 4928
rect 7114 4868 7118 4924
rect 7118 4868 7174 4924
rect 7174 4868 7178 4924
rect 7114 4864 7178 4868
rect 10822 4924 10886 4928
rect 10822 4868 10826 4924
rect 10826 4868 10882 4924
rect 10882 4868 10886 4924
rect 10822 4864 10886 4868
rect 10902 4924 10966 4928
rect 10902 4868 10906 4924
rect 10906 4868 10962 4924
rect 10962 4868 10966 4924
rect 10902 4864 10966 4868
rect 10982 4924 11046 4928
rect 10982 4868 10986 4924
rect 10986 4868 11042 4924
rect 11042 4868 11046 4924
rect 10982 4864 11046 4868
rect 11062 4924 11126 4928
rect 11062 4868 11066 4924
rect 11066 4868 11122 4924
rect 11122 4868 11126 4924
rect 11062 4864 11126 4868
rect 14770 4924 14834 4928
rect 14770 4868 14774 4924
rect 14774 4868 14830 4924
rect 14830 4868 14834 4924
rect 14770 4864 14834 4868
rect 14850 4924 14914 4928
rect 14850 4868 14854 4924
rect 14854 4868 14910 4924
rect 14910 4868 14914 4924
rect 14850 4864 14914 4868
rect 14930 4924 14994 4928
rect 14930 4868 14934 4924
rect 14934 4868 14990 4924
rect 14990 4868 14994 4924
rect 14930 4864 14994 4868
rect 15010 4924 15074 4928
rect 15010 4868 15014 4924
rect 15014 4868 15070 4924
rect 15070 4868 15074 4924
rect 15010 4864 15074 4868
rect 8708 4660 8772 4724
rect 4900 4380 4964 4384
rect 4900 4324 4904 4380
rect 4904 4324 4960 4380
rect 4960 4324 4964 4380
rect 4900 4320 4964 4324
rect 4980 4380 5044 4384
rect 4980 4324 4984 4380
rect 4984 4324 5040 4380
rect 5040 4324 5044 4380
rect 4980 4320 5044 4324
rect 5060 4380 5124 4384
rect 5060 4324 5064 4380
rect 5064 4324 5120 4380
rect 5120 4324 5124 4380
rect 5060 4320 5124 4324
rect 5140 4380 5204 4384
rect 5140 4324 5144 4380
rect 5144 4324 5200 4380
rect 5200 4324 5204 4380
rect 5140 4320 5204 4324
rect 8848 4380 8912 4384
rect 8848 4324 8852 4380
rect 8852 4324 8908 4380
rect 8908 4324 8912 4380
rect 8848 4320 8912 4324
rect 8928 4380 8992 4384
rect 8928 4324 8932 4380
rect 8932 4324 8988 4380
rect 8988 4324 8992 4380
rect 8928 4320 8992 4324
rect 9008 4380 9072 4384
rect 9008 4324 9012 4380
rect 9012 4324 9068 4380
rect 9068 4324 9072 4380
rect 9008 4320 9072 4324
rect 9088 4380 9152 4384
rect 9088 4324 9092 4380
rect 9092 4324 9148 4380
rect 9148 4324 9152 4380
rect 9088 4320 9152 4324
rect 12796 4380 12860 4384
rect 12796 4324 12800 4380
rect 12800 4324 12856 4380
rect 12856 4324 12860 4380
rect 12796 4320 12860 4324
rect 12876 4380 12940 4384
rect 12876 4324 12880 4380
rect 12880 4324 12936 4380
rect 12936 4324 12940 4380
rect 12876 4320 12940 4324
rect 12956 4380 13020 4384
rect 12956 4324 12960 4380
rect 12960 4324 13016 4380
rect 13016 4324 13020 4380
rect 12956 4320 13020 4324
rect 13036 4380 13100 4384
rect 13036 4324 13040 4380
rect 13040 4324 13096 4380
rect 13096 4324 13100 4380
rect 13036 4320 13100 4324
rect 2636 4252 2700 4316
rect 3924 4040 3988 4044
rect 5580 4116 5644 4180
rect 3924 3984 3974 4040
rect 3974 3984 3988 4040
rect 3924 3980 3988 3984
rect 8340 3980 8404 4044
rect 2926 3836 2990 3840
rect 2926 3780 2930 3836
rect 2930 3780 2986 3836
rect 2986 3780 2990 3836
rect 2926 3776 2990 3780
rect 3006 3836 3070 3840
rect 3006 3780 3010 3836
rect 3010 3780 3066 3836
rect 3066 3780 3070 3836
rect 3006 3776 3070 3780
rect 3086 3836 3150 3840
rect 3086 3780 3090 3836
rect 3090 3780 3146 3836
rect 3146 3780 3150 3836
rect 3086 3776 3150 3780
rect 3166 3836 3230 3840
rect 3166 3780 3170 3836
rect 3170 3780 3226 3836
rect 3226 3780 3230 3836
rect 3166 3776 3230 3780
rect 6874 3836 6938 3840
rect 6874 3780 6878 3836
rect 6878 3780 6934 3836
rect 6934 3780 6938 3836
rect 6874 3776 6938 3780
rect 6954 3836 7018 3840
rect 6954 3780 6958 3836
rect 6958 3780 7014 3836
rect 7014 3780 7018 3836
rect 6954 3776 7018 3780
rect 7034 3836 7098 3840
rect 7034 3780 7038 3836
rect 7038 3780 7094 3836
rect 7094 3780 7098 3836
rect 7034 3776 7098 3780
rect 7114 3836 7178 3840
rect 7114 3780 7118 3836
rect 7118 3780 7174 3836
rect 7174 3780 7178 3836
rect 7114 3776 7178 3780
rect 10822 3836 10886 3840
rect 10822 3780 10826 3836
rect 10826 3780 10882 3836
rect 10882 3780 10886 3836
rect 10822 3776 10886 3780
rect 10902 3836 10966 3840
rect 10902 3780 10906 3836
rect 10906 3780 10962 3836
rect 10962 3780 10966 3836
rect 10902 3776 10966 3780
rect 10982 3836 11046 3840
rect 10982 3780 10986 3836
rect 10986 3780 11042 3836
rect 11042 3780 11046 3836
rect 10982 3776 11046 3780
rect 11062 3836 11126 3840
rect 11062 3780 11066 3836
rect 11066 3780 11122 3836
rect 11122 3780 11126 3836
rect 11062 3776 11126 3780
rect 14770 3836 14834 3840
rect 14770 3780 14774 3836
rect 14774 3780 14830 3836
rect 14830 3780 14834 3836
rect 14770 3776 14834 3780
rect 14850 3836 14914 3840
rect 14850 3780 14854 3836
rect 14854 3780 14910 3836
rect 14910 3780 14914 3836
rect 14850 3776 14914 3780
rect 14930 3836 14994 3840
rect 14930 3780 14934 3836
rect 14934 3780 14990 3836
rect 14990 3780 14994 3836
rect 14930 3776 14994 3780
rect 15010 3836 15074 3840
rect 15010 3780 15014 3836
rect 15014 3780 15070 3836
rect 15070 3780 15074 3836
rect 15010 3776 15074 3780
rect 4108 3572 4172 3636
rect 3740 3436 3804 3500
rect 4900 3292 4964 3296
rect 4900 3236 4904 3292
rect 4904 3236 4960 3292
rect 4960 3236 4964 3292
rect 4900 3232 4964 3236
rect 4980 3292 5044 3296
rect 4980 3236 4984 3292
rect 4984 3236 5040 3292
rect 5040 3236 5044 3292
rect 4980 3232 5044 3236
rect 5060 3292 5124 3296
rect 5060 3236 5064 3292
rect 5064 3236 5120 3292
rect 5120 3236 5124 3292
rect 5060 3232 5124 3236
rect 5140 3292 5204 3296
rect 5140 3236 5144 3292
rect 5144 3236 5200 3292
rect 5200 3236 5204 3292
rect 5140 3232 5204 3236
rect 8848 3292 8912 3296
rect 8848 3236 8852 3292
rect 8852 3236 8908 3292
rect 8908 3236 8912 3292
rect 8848 3232 8912 3236
rect 8928 3292 8992 3296
rect 8928 3236 8932 3292
rect 8932 3236 8988 3292
rect 8988 3236 8992 3292
rect 8928 3232 8992 3236
rect 9008 3292 9072 3296
rect 9008 3236 9012 3292
rect 9012 3236 9068 3292
rect 9068 3236 9072 3292
rect 9008 3232 9072 3236
rect 9088 3292 9152 3296
rect 9088 3236 9092 3292
rect 9092 3236 9148 3292
rect 9148 3236 9152 3292
rect 9088 3232 9152 3236
rect 12796 3292 12860 3296
rect 12796 3236 12800 3292
rect 12800 3236 12856 3292
rect 12856 3236 12860 3292
rect 12796 3232 12860 3236
rect 12876 3292 12940 3296
rect 12876 3236 12880 3292
rect 12880 3236 12936 3292
rect 12936 3236 12940 3292
rect 12876 3232 12940 3236
rect 12956 3292 13020 3296
rect 12956 3236 12960 3292
rect 12960 3236 13016 3292
rect 13016 3236 13020 3292
rect 12956 3232 13020 3236
rect 13036 3292 13100 3296
rect 13036 3236 13040 3292
rect 13040 3236 13096 3292
rect 13096 3236 13100 3292
rect 13036 3232 13100 3236
rect 9812 3028 9876 3092
rect 2926 2748 2990 2752
rect 2926 2692 2930 2748
rect 2930 2692 2986 2748
rect 2986 2692 2990 2748
rect 2926 2688 2990 2692
rect 3006 2748 3070 2752
rect 3006 2692 3010 2748
rect 3010 2692 3066 2748
rect 3066 2692 3070 2748
rect 3006 2688 3070 2692
rect 3086 2748 3150 2752
rect 3086 2692 3090 2748
rect 3090 2692 3146 2748
rect 3146 2692 3150 2748
rect 3086 2688 3150 2692
rect 3166 2748 3230 2752
rect 3166 2692 3170 2748
rect 3170 2692 3226 2748
rect 3226 2692 3230 2748
rect 3166 2688 3230 2692
rect 6874 2748 6938 2752
rect 6874 2692 6878 2748
rect 6878 2692 6934 2748
rect 6934 2692 6938 2748
rect 6874 2688 6938 2692
rect 6954 2748 7018 2752
rect 6954 2692 6958 2748
rect 6958 2692 7014 2748
rect 7014 2692 7018 2748
rect 6954 2688 7018 2692
rect 7034 2748 7098 2752
rect 7034 2692 7038 2748
rect 7038 2692 7094 2748
rect 7094 2692 7098 2748
rect 7034 2688 7098 2692
rect 7114 2748 7178 2752
rect 7114 2692 7118 2748
rect 7118 2692 7174 2748
rect 7174 2692 7178 2748
rect 7114 2688 7178 2692
rect 10822 2748 10886 2752
rect 10822 2692 10826 2748
rect 10826 2692 10882 2748
rect 10882 2692 10886 2748
rect 10822 2688 10886 2692
rect 10902 2748 10966 2752
rect 10902 2692 10906 2748
rect 10906 2692 10962 2748
rect 10962 2692 10966 2748
rect 10902 2688 10966 2692
rect 10982 2748 11046 2752
rect 10982 2692 10986 2748
rect 10986 2692 11042 2748
rect 11042 2692 11046 2748
rect 10982 2688 11046 2692
rect 11062 2748 11126 2752
rect 11062 2692 11066 2748
rect 11066 2692 11122 2748
rect 11122 2692 11126 2748
rect 11062 2688 11126 2692
rect 14770 2748 14834 2752
rect 14770 2692 14774 2748
rect 14774 2692 14830 2748
rect 14830 2692 14834 2748
rect 14770 2688 14834 2692
rect 14850 2748 14914 2752
rect 14850 2692 14854 2748
rect 14854 2692 14910 2748
rect 14910 2692 14914 2748
rect 14850 2688 14914 2692
rect 14930 2748 14994 2752
rect 14930 2692 14934 2748
rect 14934 2692 14990 2748
rect 14990 2692 14994 2748
rect 14930 2688 14994 2692
rect 15010 2748 15074 2752
rect 15010 2692 15014 2748
rect 15014 2692 15070 2748
rect 15070 2692 15074 2748
rect 15010 2688 15074 2692
rect 4900 2204 4964 2208
rect 4900 2148 4904 2204
rect 4904 2148 4960 2204
rect 4960 2148 4964 2204
rect 4900 2144 4964 2148
rect 4980 2204 5044 2208
rect 4980 2148 4984 2204
rect 4984 2148 5040 2204
rect 5040 2148 5044 2204
rect 4980 2144 5044 2148
rect 5060 2204 5124 2208
rect 5060 2148 5064 2204
rect 5064 2148 5120 2204
rect 5120 2148 5124 2204
rect 5060 2144 5124 2148
rect 5140 2204 5204 2208
rect 5140 2148 5144 2204
rect 5144 2148 5200 2204
rect 5200 2148 5204 2204
rect 5140 2144 5204 2148
rect 8848 2204 8912 2208
rect 8848 2148 8852 2204
rect 8852 2148 8908 2204
rect 8908 2148 8912 2204
rect 8848 2144 8912 2148
rect 8928 2204 8992 2208
rect 8928 2148 8932 2204
rect 8932 2148 8988 2204
rect 8988 2148 8992 2204
rect 8928 2144 8992 2148
rect 9008 2204 9072 2208
rect 9008 2148 9012 2204
rect 9012 2148 9068 2204
rect 9068 2148 9072 2204
rect 9008 2144 9072 2148
rect 9088 2204 9152 2208
rect 9088 2148 9092 2204
rect 9092 2148 9148 2204
rect 9148 2148 9152 2204
rect 9088 2144 9152 2148
rect 12796 2204 12860 2208
rect 12796 2148 12800 2204
rect 12800 2148 12856 2204
rect 12856 2148 12860 2204
rect 12796 2144 12860 2148
rect 12876 2204 12940 2208
rect 12876 2148 12880 2204
rect 12880 2148 12936 2204
rect 12936 2148 12940 2204
rect 12876 2144 12940 2148
rect 12956 2204 13020 2208
rect 12956 2148 12960 2204
rect 12960 2148 13016 2204
rect 13016 2148 13020 2204
rect 12956 2144 13020 2148
rect 13036 2204 13100 2208
rect 13036 2148 13040 2204
rect 13040 2148 13096 2204
rect 13096 2148 13100 2204
rect 13036 2144 13100 2148
rect 2926 1660 2990 1664
rect 2926 1604 2930 1660
rect 2930 1604 2986 1660
rect 2986 1604 2990 1660
rect 2926 1600 2990 1604
rect 3006 1660 3070 1664
rect 3006 1604 3010 1660
rect 3010 1604 3066 1660
rect 3066 1604 3070 1660
rect 3006 1600 3070 1604
rect 3086 1660 3150 1664
rect 3086 1604 3090 1660
rect 3090 1604 3146 1660
rect 3146 1604 3150 1660
rect 3086 1600 3150 1604
rect 3166 1660 3230 1664
rect 3166 1604 3170 1660
rect 3170 1604 3226 1660
rect 3226 1604 3230 1660
rect 3166 1600 3230 1604
rect 6874 1660 6938 1664
rect 6874 1604 6878 1660
rect 6878 1604 6934 1660
rect 6934 1604 6938 1660
rect 6874 1600 6938 1604
rect 6954 1660 7018 1664
rect 6954 1604 6958 1660
rect 6958 1604 7014 1660
rect 7014 1604 7018 1660
rect 6954 1600 7018 1604
rect 7034 1660 7098 1664
rect 7034 1604 7038 1660
rect 7038 1604 7094 1660
rect 7094 1604 7098 1660
rect 7034 1600 7098 1604
rect 7114 1660 7178 1664
rect 7114 1604 7118 1660
rect 7118 1604 7174 1660
rect 7174 1604 7178 1660
rect 7114 1600 7178 1604
rect 10822 1660 10886 1664
rect 10822 1604 10826 1660
rect 10826 1604 10882 1660
rect 10882 1604 10886 1660
rect 10822 1600 10886 1604
rect 10902 1660 10966 1664
rect 10902 1604 10906 1660
rect 10906 1604 10962 1660
rect 10962 1604 10966 1660
rect 10902 1600 10966 1604
rect 10982 1660 11046 1664
rect 10982 1604 10986 1660
rect 10986 1604 11042 1660
rect 11042 1604 11046 1660
rect 10982 1600 11046 1604
rect 11062 1660 11126 1664
rect 11062 1604 11066 1660
rect 11066 1604 11122 1660
rect 11122 1604 11126 1660
rect 11062 1600 11126 1604
rect 14770 1660 14834 1664
rect 14770 1604 14774 1660
rect 14774 1604 14830 1660
rect 14830 1604 14834 1660
rect 14770 1600 14834 1604
rect 14850 1660 14914 1664
rect 14850 1604 14854 1660
rect 14854 1604 14910 1660
rect 14910 1604 14914 1660
rect 14850 1600 14914 1604
rect 14930 1660 14994 1664
rect 14930 1604 14934 1660
rect 14934 1604 14990 1660
rect 14990 1604 14994 1660
rect 14930 1600 14994 1604
rect 15010 1660 15074 1664
rect 15010 1604 15014 1660
rect 15014 1604 15070 1660
rect 15070 1604 15074 1660
rect 15010 1600 15074 1604
rect 4900 1116 4964 1120
rect 4900 1060 4904 1116
rect 4904 1060 4960 1116
rect 4960 1060 4964 1116
rect 4900 1056 4964 1060
rect 4980 1116 5044 1120
rect 4980 1060 4984 1116
rect 4984 1060 5040 1116
rect 5040 1060 5044 1116
rect 4980 1056 5044 1060
rect 5060 1116 5124 1120
rect 5060 1060 5064 1116
rect 5064 1060 5120 1116
rect 5120 1060 5124 1116
rect 5060 1056 5124 1060
rect 5140 1116 5204 1120
rect 5140 1060 5144 1116
rect 5144 1060 5200 1116
rect 5200 1060 5204 1116
rect 5140 1056 5204 1060
rect 8848 1116 8912 1120
rect 8848 1060 8852 1116
rect 8852 1060 8908 1116
rect 8908 1060 8912 1116
rect 8848 1056 8912 1060
rect 8928 1116 8992 1120
rect 8928 1060 8932 1116
rect 8932 1060 8988 1116
rect 8988 1060 8992 1116
rect 8928 1056 8992 1060
rect 9008 1116 9072 1120
rect 9008 1060 9012 1116
rect 9012 1060 9068 1116
rect 9068 1060 9072 1116
rect 9008 1056 9072 1060
rect 9088 1116 9152 1120
rect 9088 1060 9092 1116
rect 9092 1060 9148 1116
rect 9148 1060 9152 1116
rect 9088 1056 9152 1060
rect 12796 1116 12860 1120
rect 12796 1060 12800 1116
rect 12800 1060 12856 1116
rect 12856 1060 12860 1116
rect 12796 1056 12860 1060
rect 12876 1116 12940 1120
rect 12876 1060 12880 1116
rect 12880 1060 12936 1116
rect 12936 1060 12940 1116
rect 12876 1056 12940 1060
rect 12956 1116 13020 1120
rect 12956 1060 12960 1116
rect 12960 1060 13016 1116
rect 13016 1060 13020 1116
rect 12956 1056 13020 1060
rect 13036 1116 13100 1120
rect 13036 1060 13040 1116
rect 13040 1060 13096 1116
rect 13096 1060 13100 1116
rect 13036 1056 13100 1060
<< metal4 >>
rect 2918 22336 3238 22896
rect 2918 22272 2926 22336
rect 2990 22272 3006 22336
rect 3070 22272 3086 22336
rect 3150 22272 3166 22336
rect 3230 22272 3238 22336
rect 2918 21248 3238 22272
rect 2918 21184 2926 21248
rect 2990 21184 3006 21248
rect 3070 21184 3086 21248
rect 3150 21184 3166 21248
rect 3230 21184 3238 21248
rect 2918 20160 3238 21184
rect 2918 20096 2926 20160
rect 2990 20096 3006 20160
rect 3070 20096 3086 20160
rect 3150 20096 3166 20160
rect 3230 20096 3238 20160
rect 2918 19072 3238 20096
rect 2918 19008 2926 19072
rect 2990 19008 3006 19072
rect 3070 19008 3086 19072
rect 3150 19008 3166 19072
rect 3230 19008 3238 19072
rect 2918 17984 3238 19008
rect 2918 17920 2926 17984
rect 2990 17920 3006 17984
rect 3070 17920 3086 17984
rect 3150 17920 3166 17984
rect 3230 17920 3238 17984
rect 2918 16896 3238 17920
rect 2918 16832 2926 16896
rect 2990 16832 3006 16896
rect 3070 16832 3086 16896
rect 3150 16832 3166 16896
rect 3230 16832 3238 16896
rect 2918 15808 3238 16832
rect 2918 15744 2926 15808
rect 2990 15744 3006 15808
rect 3070 15744 3086 15808
rect 3150 15744 3166 15808
rect 3230 15744 3238 15808
rect 2918 14720 3238 15744
rect 2918 14656 2926 14720
rect 2990 14656 3006 14720
rect 3070 14656 3086 14720
rect 3150 14656 3166 14720
rect 3230 14656 3238 14720
rect 2918 13632 3238 14656
rect 4892 22880 5212 22896
rect 4892 22816 4900 22880
rect 4964 22816 4980 22880
rect 5044 22816 5060 22880
rect 5124 22816 5140 22880
rect 5204 22816 5212 22880
rect 4892 21792 5212 22816
rect 4892 21728 4900 21792
rect 4964 21728 4980 21792
rect 5044 21728 5060 21792
rect 5124 21728 5140 21792
rect 5204 21728 5212 21792
rect 4892 20704 5212 21728
rect 4892 20640 4900 20704
rect 4964 20640 4980 20704
rect 5044 20640 5060 20704
rect 5124 20640 5140 20704
rect 5204 20640 5212 20704
rect 4892 19616 5212 20640
rect 4892 19552 4900 19616
rect 4964 19552 4980 19616
rect 5044 19552 5060 19616
rect 5124 19552 5140 19616
rect 5204 19552 5212 19616
rect 4892 18528 5212 19552
rect 4892 18464 4900 18528
rect 4964 18464 4980 18528
rect 5044 18464 5060 18528
rect 5124 18464 5140 18528
rect 5204 18464 5212 18528
rect 4892 17440 5212 18464
rect 4892 17376 4900 17440
rect 4964 17376 4980 17440
rect 5044 17376 5060 17440
rect 5124 17376 5140 17440
rect 5204 17376 5212 17440
rect 4892 16352 5212 17376
rect 4892 16288 4900 16352
rect 4964 16288 4980 16352
rect 5044 16288 5060 16352
rect 5124 16288 5140 16352
rect 5204 16288 5212 16352
rect 4892 15264 5212 16288
rect 6866 22336 7186 22896
rect 6866 22272 6874 22336
rect 6938 22272 6954 22336
rect 7018 22272 7034 22336
rect 7098 22272 7114 22336
rect 7178 22272 7186 22336
rect 6866 21248 7186 22272
rect 6866 21184 6874 21248
rect 6938 21184 6954 21248
rect 7018 21184 7034 21248
rect 7098 21184 7114 21248
rect 7178 21184 7186 21248
rect 6866 20160 7186 21184
rect 6866 20096 6874 20160
rect 6938 20096 6954 20160
rect 7018 20096 7034 20160
rect 7098 20096 7114 20160
rect 7178 20096 7186 20160
rect 6866 19072 7186 20096
rect 6866 19008 6874 19072
rect 6938 19008 6954 19072
rect 7018 19008 7034 19072
rect 7098 19008 7114 19072
rect 7178 19008 7186 19072
rect 6866 17984 7186 19008
rect 6866 17920 6874 17984
rect 6938 17920 6954 17984
rect 7018 17920 7034 17984
rect 7098 17920 7114 17984
rect 7178 17920 7186 17984
rect 6866 16896 7186 17920
rect 6866 16832 6874 16896
rect 6938 16832 6954 16896
rect 7018 16832 7034 16896
rect 7098 16832 7114 16896
rect 7178 16832 7186 16896
rect 6866 15808 7186 16832
rect 6866 15744 6874 15808
rect 6938 15744 6954 15808
rect 7018 15744 7034 15808
rect 7098 15744 7114 15808
rect 7178 15744 7186 15808
rect 5395 15468 5461 15469
rect 5395 15404 5396 15468
rect 5460 15404 5461 15468
rect 5395 15403 5461 15404
rect 6499 15468 6565 15469
rect 6499 15404 6500 15468
rect 6564 15404 6565 15468
rect 6499 15403 6565 15404
rect 4892 15200 4900 15264
rect 4964 15200 4980 15264
rect 5044 15200 5060 15264
rect 5124 15200 5140 15264
rect 5204 15200 5212 15264
rect 3923 14380 3989 14381
rect 3923 14316 3924 14380
rect 3988 14316 3989 14380
rect 3923 14315 3989 14316
rect 2918 13568 2926 13632
rect 2990 13568 3006 13632
rect 3070 13568 3086 13632
rect 3150 13568 3166 13632
rect 3230 13568 3238 13632
rect 2918 12544 3238 13568
rect 2918 12480 2926 12544
rect 2990 12480 3006 12544
rect 3070 12480 3086 12544
rect 3150 12480 3166 12544
rect 3230 12480 3238 12544
rect 2918 11456 3238 12480
rect 3555 11796 3621 11797
rect 3555 11732 3556 11796
rect 3620 11732 3621 11796
rect 3555 11731 3621 11732
rect 2918 11392 2926 11456
rect 2990 11392 3006 11456
rect 3070 11392 3086 11456
rect 3150 11392 3166 11456
rect 3230 11392 3238 11456
rect 2635 11116 2701 11117
rect 2635 11052 2636 11116
rect 2700 11052 2701 11116
rect 2635 11051 2701 11052
rect 2638 10029 2698 11051
rect 2918 10368 3238 11392
rect 2918 10304 2926 10368
rect 2990 10304 3006 10368
rect 3070 10304 3086 10368
rect 3150 10304 3166 10368
rect 3230 10304 3238 10368
rect 2635 10028 2701 10029
rect 2635 9964 2636 10028
rect 2700 9964 2701 10028
rect 2635 9963 2701 9964
rect 2638 4317 2698 9963
rect 2918 9280 3238 10304
rect 2918 9216 2926 9280
rect 2990 9216 3006 9280
rect 3070 9216 3086 9280
rect 3150 9216 3166 9280
rect 3230 9216 3238 9280
rect 2918 8192 3238 9216
rect 2918 8128 2926 8192
rect 2990 8128 3006 8192
rect 3070 8128 3086 8192
rect 3150 8128 3166 8192
rect 3230 8128 3238 8192
rect 2918 7104 3238 8128
rect 2918 7040 2926 7104
rect 2990 7040 3006 7104
rect 3070 7040 3086 7104
rect 3150 7040 3166 7104
rect 3230 7040 3238 7104
rect 2918 6016 3238 7040
rect 2918 5952 2926 6016
rect 2990 5952 3006 6016
rect 3070 5952 3086 6016
rect 3150 5952 3166 6016
rect 3230 5952 3238 6016
rect 2918 4928 3238 5952
rect 3558 5405 3618 11731
rect 3739 11524 3805 11525
rect 3739 11460 3740 11524
rect 3804 11460 3805 11524
rect 3739 11459 3805 11460
rect 3555 5404 3621 5405
rect 3555 5340 3556 5404
rect 3620 5340 3621 5404
rect 3555 5339 3621 5340
rect 2918 4864 2926 4928
rect 2990 4864 3006 4928
rect 3070 4864 3086 4928
rect 3150 4864 3166 4928
rect 3230 4864 3238 4928
rect 2635 4316 2701 4317
rect 2635 4252 2636 4316
rect 2700 4252 2701 4316
rect 2635 4251 2701 4252
rect 2918 3840 3238 4864
rect 2918 3776 2926 3840
rect 2990 3776 3006 3840
rect 3070 3776 3086 3840
rect 3150 3776 3166 3840
rect 3230 3776 3238 3840
rect 2918 2752 3238 3776
rect 3742 3501 3802 11459
rect 3926 4045 3986 14315
rect 4892 14176 5212 15200
rect 4892 14112 4900 14176
rect 4964 14112 4980 14176
rect 5044 14112 5060 14176
rect 5124 14112 5140 14176
rect 5204 14112 5212 14176
rect 4892 13088 5212 14112
rect 4892 13024 4900 13088
rect 4964 13024 4980 13088
rect 5044 13024 5060 13088
rect 5124 13024 5140 13088
rect 5204 13024 5212 13088
rect 4892 12000 5212 13024
rect 4892 11936 4900 12000
rect 4964 11936 4980 12000
rect 5044 11936 5060 12000
rect 5124 11936 5140 12000
rect 5204 11936 5212 12000
rect 4892 10912 5212 11936
rect 4892 10848 4900 10912
rect 4964 10848 4980 10912
rect 5044 10848 5060 10912
rect 5124 10848 5140 10912
rect 5204 10848 5212 10912
rect 4892 9824 5212 10848
rect 4892 9760 4900 9824
rect 4964 9760 4980 9824
rect 5044 9760 5060 9824
rect 5124 9760 5140 9824
rect 5204 9760 5212 9824
rect 4659 9620 4725 9621
rect 4659 9556 4660 9620
rect 4724 9556 4725 9620
rect 4659 9555 4725 9556
rect 4107 7036 4173 7037
rect 4107 6972 4108 7036
rect 4172 6972 4173 7036
rect 4107 6971 4173 6972
rect 3923 4044 3989 4045
rect 3923 3980 3924 4044
rect 3988 3980 3989 4044
rect 3923 3979 3989 3980
rect 4110 3637 4170 6971
rect 4662 4997 4722 9555
rect 4892 8736 5212 9760
rect 4892 8672 4900 8736
rect 4964 8672 4980 8736
rect 5044 8672 5060 8736
rect 5124 8672 5140 8736
rect 5204 8672 5212 8736
rect 4892 7648 5212 8672
rect 4892 7584 4900 7648
rect 4964 7584 4980 7648
rect 5044 7584 5060 7648
rect 5124 7584 5140 7648
rect 5204 7584 5212 7648
rect 4892 6560 5212 7584
rect 4892 6496 4900 6560
rect 4964 6496 4980 6560
rect 5044 6496 5060 6560
rect 5124 6496 5140 6560
rect 5204 6496 5212 6560
rect 4892 5472 5212 6496
rect 4892 5408 4900 5472
rect 4964 5408 4980 5472
rect 5044 5408 5060 5472
rect 5124 5408 5140 5472
rect 5204 5408 5212 5472
rect 4659 4996 4725 4997
rect 4659 4932 4660 4996
rect 4724 4932 4725 4996
rect 4659 4931 4725 4932
rect 4892 4384 5212 5408
rect 5398 5405 5458 15403
rect 5947 11116 6013 11117
rect 5947 11052 5948 11116
rect 6012 11052 6013 11116
rect 5947 11051 6013 11052
rect 5579 8396 5645 8397
rect 5579 8332 5580 8396
rect 5644 8332 5645 8396
rect 5579 8331 5645 8332
rect 5395 5404 5461 5405
rect 5395 5340 5396 5404
rect 5460 5340 5461 5404
rect 5395 5339 5461 5340
rect 4892 4320 4900 4384
rect 4964 4320 4980 4384
rect 5044 4320 5060 4384
rect 5124 4320 5140 4384
rect 5204 4320 5212 4384
rect 4107 3636 4173 3637
rect 4107 3572 4108 3636
rect 4172 3572 4173 3636
rect 4107 3571 4173 3572
rect 3739 3500 3805 3501
rect 3739 3436 3740 3500
rect 3804 3436 3805 3500
rect 3739 3435 3805 3436
rect 2918 2688 2926 2752
rect 2990 2688 3006 2752
rect 3070 2688 3086 2752
rect 3150 2688 3166 2752
rect 3230 2688 3238 2752
rect 2918 1664 3238 2688
rect 2918 1600 2926 1664
rect 2990 1600 3006 1664
rect 3070 1600 3086 1664
rect 3150 1600 3166 1664
rect 3230 1600 3238 1664
rect 2918 1040 3238 1600
rect 4892 3296 5212 4320
rect 5582 4181 5642 8331
rect 5763 8124 5829 8125
rect 5763 8060 5764 8124
rect 5828 8060 5829 8124
rect 5763 8059 5829 8060
rect 5766 6629 5826 8059
rect 5950 7581 6010 11051
rect 6131 8124 6197 8125
rect 6131 8060 6132 8124
rect 6196 8060 6197 8124
rect 6131 8059 6197 8060
rect 6315 8124 6381 8125
rect 6315 8060 6316 8124
rect 6380 8060 6381 8124
rect 6315 8059 6381 8060
rect 5947 7580 6013 7581
rect 5947 7516 5948 7580
rect 6012 7516 6013 7580
rect 5947 7515 6013 7516
rect 6134 7173 6194 8059
rect 6131 7172 6197 7173
rect 6131 7108 6132 7172
rect 6196 7108 6197 7172
rect 6131 7107 6197 7108
rect 6318 6901 6378 8059
rect 6502 7173 6562 15403
rect 6866 14720 7186 15744
rect 8840 22880 9160 22896
rect 8840 22816 8848 22880
rect 8912 22816 8928 22880
rect 8992 22816 9008 22880
rect 9072 22816 9088 22880
rect 9152 22816 9160 22880
rect 8840 21792 9160 22816
rect 8840 21728 8848 21792
rect 8912 21728 8928 21792
rect 8992 21728 9008 21792
rect 9072 21728 9088 21792
rect 9152 21728 9160 21792
rect 8840 20704 9160 21728
rect 8840 20640 8848 20704
rect 8912 20640 8928 20704
rect 8992 20640 9008 20704
rect 9072 20640 9088 20704
rect 9152 20640 9160 20704
rect 8840 19616 9160 20640
rect 8840 19552 8848 19616
rect 8912 19552 8928 19616
rect 8992 19552 9008 19616
rect 9072 19552 9088 19616
rect 9152 19552 9160 19616
rect 8840 18528 9160 19552
rect 8840 18464 8848 18528
rect 8912 18464 8928 18528
rect 8992 18464 9008 18528
rect 9072 18464 9088 18528
rect 9152 18464 9160 18528
rect 8840 17440 9160 18464
rect 8840 17376 8848 17440
rect 8912 17376 8928 17440
rect 8992 17376 9008 17440
rect 9072 17376 9088 17440
rect 9152 17376 9160 17440
rect 8840 16352 9160 17376
rect 8840 16288 8848 16352
rect 8912 16288 8928 16352
rect 8992 16288 9008 16352
rect 9072 16288 9088 16352
rect 9152 16288 9160 16352
rect 8840 15264 9160 16288
rect 8840 15200 8848 15264
rect 8912 15200 8928 15264
rect 8992 15200 9008 15264
rect 9072 15200 9088 15264
rect 9152 15200 9160 15264
rect 7419 14924 7485 14925
rect 7419 14860 7420 14924
rect 7484 14860 7485 14924
rect 7419 14859 7485 14860
rect 6866 14656 6874 14720
rect 6938 14656 6954 14720
rect 7018 14656 7034 14720
rect 7098 14656 7114 14720
rect 7178 14656 7186 14720
rect 6866 13632 7186 14656
rect 6866 13568 6874 13632
rect 6938 13568 6954 13632
rect 7018 13568 7034 13632
rect 7098 13568 7114 13632
rect 7178 13568 7186 13632
rect 6866 12544 7186 13568
rect 6866 12480 6874 12544
rect 6938 12480 6954 12544
rect 7018 12480 7034 12544
rect 7098 12480 7114 12544
rect 7178 12480 7186 12544
rect 6866 11456 7186 12480
rect 6866 11392 6874 11456
rect 6938 11392 6954 11456
rect 7018 11392 7034 11456
rect 7098 11392 7114 11456
rect 7178 11392 7186 11456
rect 6866 10368 7186 11392
rect 6866 10304 6874 10368
rect 6938 10304 6954 10368
rect 7018 10304 7034 10368
rect 7098 10304 7114 10368
rect 7178 10304 7186 10368
rect 6866 9280 7186 10304
rect 7422 10301 7482 14859
rect 8840 14176 9160 15200
rect 8840 14112 8848 14176
rect 8912 14112 8928 14176
rect 8992 14112 9008 14176
rect 9072 14112 9088 14176
rect 9152 14112 9160 14176
rect 8707 13428 8773 13429
rect 8707 13364 8708 13428
rect 8772 13364 8773 13428
rect 8707 13363 8773 13364
rect 8523 12068 8589 12069
rect 8523 12004 8524 12068
rect 8588 12004 8589 12068
rect 8523 12003 8589 12004
rect 8155 10708 8221 10709
rect 8155 10644 8156 10708
rect 8220 10644 8221 10708
rect 8155 10643 8221 10644
rect 7971 10436 8037 10437
rect 7971 10372 7972 10436
rect 8036 10372 8037 10436
rect 7971 10371 8037 10372
rect 7419 10300 7485 10301
rect 7419 10236 7420 10300
rect 7484 10236 7485 10300
rect 7419 10235 7485 10236
rect 6866 9216 6874 9280
rect 6938 9216 6954 9280
rect 7018 9216 7034 9280
rect 7098 9216 7114 9280
rect 7178 9216 7186 9280
rect 6683 8804 6749 8805
rect 6683 8740 6684 8804
rect 6748 8740 6749 8804
rect 6683 8739 6749 8740
rect 6499 7172 6565 7173
rect 6499 7108 6500 7172
rect 6564 7108 6565 7172
rect 6499 7107 6565 7108
rect 6315 6900 6381 6901
rect 6315 6836 6316 6900
rect 6380 6836 6381 6900
rect 6315 6835 6381 6836
rect 5763 6628 5829 6629
rect 5763 6564 5764 6628
rect 5828 6564 5829 6628
rect 5763 6563 5829 6564
rect 6686 6493 6746 8739
rect 6866 8192 7186 9216
rect 7419 8396 7485 8397
rect 7419 8332 7420 8396
rect 7484 8332 7485 8396
rect 7419 8331 7485 8332
rect 6866 8128 6874 8192
rect 6938 8128 6954 8192
rect 7018 8128 7034 8192
rect 7098 8128 7114 8192
rect 7178 8128 7186 8192
rect 6866 7104 7186 8128
rect 6866 7040 6874 7104
rect 6938 7040 6954 7104
rect 7018 7040 7034 7104
rect 7098 7040 7114 7104
rect 7178 7040 7186 7104
rect 6683 6492 6749 6493
rect 6683 6428 6684 6492
rect 6748 6428 6749 6492
rect 6683 6427 6749 6428
rect 6866 6016 7186 7040
rect 6866 5952 6874 6016
rect 6938 5952 6954 6016
rect 7018 5952 7034 6016
rect 7098 5952 7114 6016
rect 7178 5952 7186 6016
rect 6866 4928 7186 5952
rect 7422 5269 7482 8331
rect 7974 6493 8034 10371
rect 8158 6629 8218 10643
rect 8339 8940 8405 8941
rect 8339 8876 8340 8940
rect 8404 8876 8405 8940
rect 8339 8875 8405 8876
rect 8155 6628 8221 6629
rect 8155 6564 8156 6628
rect 8220 6564 8221 6628
rect 8155 6563 8221 6564
rect 7971 6492 8037 6493
rect 7971 6428 7972 6492
rect 8036 6428 8037 6492
rect 7971 6427 8037 6428
rect 7419 5268 7485 5269
rect 7419 5204 7420 5268
rect 7484 5204 7485 5268
rect 7419 5203 7485 5204
rect 6866 4864 6874 4928
rect 6938 4864 6954 4928
rect 7018 4864 7034 4928
rect 7098 4864 7114 4928
rect 7178 4864 7186 4928
rect 5579 4180 5645 4181
rect 5579 4116 5580 4180
rect 5644 4116 5645 4180
rect 5579 4115 5645 4116
rect 4892 3232 4900 3296
rect 4964 3232 4980 3296
rect 5044 3232 5060 3296
rect 5124 3232 5140 3296
rect 5204 3232 5212 3296
rect 4892 2208 5212 3232
rect 4892 2144 4900 2208
rect 4964 2144 4980 2208
rect 5044 2144 5060 2208
rect 5124 2144 5140 2208
rect 5204 2144 5212 2208
rect 4892 1120 5212 2144
rect 4892 1056 4900 1120
rect 4964 1056 4980 1120
rect 5044 1056 5060 1120
rect 5124 1056 5140 1120
rect 5204 1056 5212 1120
rect 4892 1040 5212 1056
rect 6866 3840 7186 4864
rect 8342 4045 8402 8875
rect 8526 5405 8586 12003
rect 8710 11797 8770 13363
rect 8840 13088 9160 14112
rect 8840 13024 8848 13088
rect 8912 13024 8928 13088
rect 8992 13024 9008 13088
rect 9072 13024 9088 13088
rect 9152 13024 9160 13088
rect 8840 12000 9160 13024
rect 10814 22336 11134 22896
rect 10814 22272 10822 22336
rect 10886 22272 10902 22336
rect 10966 22272 10982 22336
rect 11046 22272 11062 22336
rect 11126 22272 11134 22336
rect 10814 21248 11134 22272
rect 10814 21184 10822 21248
rect 10886 21184 10902 21248
rect 10966 21184 10982 21248
rect 11046 21184 11062 21248
rect 11126 21184 11134 21248
rect 10814 20160 11134 21184
rect 10814 20096 10822 20160
rect 10886 20096 10902 20160
rect 10966 20096 10982 20160
rect 11046 20096 11062 20160
rect 11126 20096 11134 20160
rect 10814 19072 11134 20096
rect 10814 19008 10822 19072
rect 10886 19008 10902 19072
rect 10966 19008 10982 19072
rect 11046 19008 11062 19072
rect 11126 19008 11134 19072
rect 10814 17984 11134 19008
rect 10814 17920 10822 17984
rect 10886 17920 10902 17984
rect 10966 17920 10982 17984
rect 11046 17920 11062 17984
rect 11126 17920 11134 17984
rect 10814 16896 11134 17920
rect 10814 16832 10822 16896
rect 10886 16832 10902 16896
rect 10966 16832 10982 16896
rect 11046 16832 11062 16896
rect 11126 16832 11134 16896
rect 10814 15808 11134 16832
rect 10814 15744 10822 15808
rect 10886 15744 10902 15808
rect 10966 15744 10982 15808
rect 11046 15744 11062 15808
rect 11126 15744 11134 15808
rect 10814 14720 11134 15744
rect 10814 14656 10822 14720
rect 10886 14656 10902 14720
rect 10966 14656 10982 14720
rect 11046 14656 11062 14720
rect 11126 14656 11134 14720
rect 10814 13632 11134 14656
rect 10814 13568 10822 13632
rect 10886 13568 10902 13632
rect 10966 13568 10982 13632
rect 11046 13568 11062 13632
rect 11126 13568 11134 13632
rect 10814 12544 11134 13568
rect 10814 12480 10822 12544
rect 10886 12480 10902 12544
rect 10966 12480 10982 12544
rect 11046 12480 11062 12544
rect 11126 12480 11134 12544
rect 9259 12476 9325 12477
rect 9259 12412 9260 12476
rect 9324 12412 9325 12476
rect 9259 12411 9325 12412
rect 9443 12476 9509 12477
rect 9443 12412 9444 12476
rect 9508 12412 9509 12476
rect 9443 12411 9509 12412
rect 9262 12069 9322 12411
rect 9259 12068 9325 12069
rect 9259 12004 9260 12068
rect 9324 12004 9325 12068
rect 9259 12003 9325 12004
rect 8840 11936 8848 12000
rect 8912 11936 8928 12000
rect 8992 11936 9008 12000
rect 9072 11936 9088 12000
rect 9152 11936 9160 12000
rect 8707 11796 8773 11797
rect 8707 11732 8708 11796
rect 8772 11732 8773 11796
rect 8707 11731 8773 11732
rect 8840 10912 9160 11936
rect 8840 10848 8848 10912
rect 8912 10848 8928 10912
rect 8992 10848 9008 10912
rect 9072 10848 9088 10912
rect 9152 10848 9160 10912
rect 8840 9824 9160 10848
rect 8840 9760 8848 9824
rect 8912 9760 8928 9824
rect 8992 9760 9008 9824
rect 9072 9760 9088 9824
rect 9152 9760 9160 9824
rect 8840 8736 9160 9760
rect 9259 9212 9325 9213
rect 9259 9148 9260 9212
rect 9324 9148 9325 9212
rect 9259 9147 9325 9148
rect 8840 8672 8848 8736
rect 8912 8672 8928 8736
rect 8992 8672 9008 8736
rect 9072 8672 9088 8736
rect 9152 8672 9160 8736
rect 8707 8396 8773 8397
rect 8707 8332 8708 8396
rect 8772 8332 8773 8396
rect 8707 8331 8773 8332
rect 8523 5404 8589 5405
rect 8523 5340 8524 5404
rect 8588 5340 8589 5404
rect 8523 5339 8589 5340
rect 8710 4725 8770 8331
rect 8840 7648 9160 8672
rect 9262 8669 9322 9147
rect 9446 8805 9506 12411
rect 9811 12340 9877 12341
rect 9811 12276 9812 12340
rect 9876 12276 9877 12340
rect 9811 12275 9877 12276
rect 9814 10845 9874 12275
rect 10547 11796 10613 11797
rect 10547 11732 10548 11796
rect 10612 11732 10613 11796
rect 10547 11731 10613 11732
rect 9811 10844 9877 10845
rect 9811 10780 9812 10844
rect 9876 10780 9877 10844
rect 9811 10779 9877 10780
rect 9627 9756 9693 9757
rect 9627 9692 9628 9756
rect 9692 9692 9693 9756
rect 9627 9691 9693 9692
rect 9443 8804 9509 8805
rect 9443 8740 9444 8804
rect 9508 8740 9509 8804
rect 9443 8739 9509 8740
rect 9259 8668 9325 8669
rect 9259 8604 9260 8668
rect 9324 8604 9325 8668
rect 9259 8603 9325 8604
rect 9446 8397 9506 8739
rect 9443 8396 9509 8397
rect 9443 8332 9444 8396
rect 9508 8332 9509 8396
rect 9443 8331 9509 8332
rect 8840 7584 8848 7648
rect 8912 7584 8928 7648
rect 8992 7584 9008 7648
rect 9072 7584 9088 7648
rect 9152 7584 9160 7648
rect 8840 6560 9160 7584
rect 8840 6496 8848 6560
rect 8912 6496 8928 6560
rect 8992 6496 9008 6560
rect 9072 6496 9088 6560
rect 9152 6496 9160 6560
rect 8840 5472 9160 6496
rect 9630 5813 9690 9691
rect 9995 9484 10061 9485
rect 9995 9420 9996 9484
rect 10060 9420 10061 9484
rect 9995 9419 10061 9420
rect 9811 8396 9877 8397
rect 9811 8332 9812 8396
rect 9876 8332 9877 8396
rect 9811 8331 9877 8332
rect 9627 5812 9693 5813
rect 9627 5748 9628 5812
rect 9692 5748 9693 5812
rect 9627 5747 9693 5748
rect 8840 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9008 5472
rect 9072 5408 9088 5472
rect 9152 5408 9160 5472
rect 8707 4724 8773 4725
rect 8707 4660 8708 4724
rect 8772 4660 8773 4724
rect 8707 4659 8773 4660
rect 8840 4384 9160 5408
rect 8840 4320 8848 4384
rect 8912 4320 8928 4384
rect 8992 4320 9008 4384
rect 9072 4320 9088 4384
rect 9152 4320 9160 4384
rect 8339 4044 8405 4045
rect 8339 3980 8340 4044
rect 8404 3980 8405 4044
rect 8339 3979 8405 3980
rect 6866 3776 6874 3840
rect 6938 3776 6954 3840
rect 7018 3776 7034 3840
rect 7098 3776 7114 3840
rect 7178 3776 7186 3840
rect 6866 2752 7186 3776
rect 6866 2688 6874 2752
rect 6938 2688 6954 2752
rect 7018 2688 7034 2752
rect 7098 2688 7114 2752
rect 7178 2688 7186 2752
rect 6866 1664 7186 2688
rect 6866 1600 6874 1664
rect 6938 1600 6954 1664
rect 7018 1600 7034 1664
rect 7098 1600 7114 1664
rect 7178 1600 7186 1664
rect 6866 1040 7186 1600
rect 8840 3296 9160 4320
rect 8840 3232 8848 3296
rect 8912 3232 8928 3296
rect 8992 3232 9008 3296
rect 9072 3232 9088 3296
rect 9152 3232 9160 3296
rect 8840 2208 9160 3232
rect 9814 3093 9874 8331
rect 9998 7581 10058 9419
rect 10179 9212 10245 9213
rect 10179 9148 10180 9212
rect 10244 9148 10245 9212
rect 10179 9147 10245 9148
rect 10363 9212 10429 9213
rect 10363 9148 10364 9212
rect 10428 9148 10429 9212
rect 10363 9147 10429 9148
rect 10182 7717 10242 9147
rect 10366 7853 10426 9147
rect 10550 8125 10610 11731
rect 10814 11456 11134 12480
rect 10814 11392 10822 11456
rect 10886 11392 10902 11456
rect 10966 11392 10982 11456
rect 11046 11392 11062 11456
rect 11126 11392 11134 11456
rect 10814 10368 11134 11392
rect 10814 10304 10822 10368
rect 10886 10304 10902 10368
rect 10966 10304 10982 10368
rect 11046 10304 11062 10368
rect 11126 10304 11134 10368
rect 10814 9280 11134 10304
rect 10814 9216 10822 9280
rect 10886 9216 10902 9280
rect 10966 9216 10982 9280
rect 11046 9216 11062 9280
rect 11126 9216 11134 9280
rect 10814 8192 11134 9216
rect 12788 22880 13108 22896
rect 12788 22816 12796 22880
rect 12860 22816 12876 22880
rect 12940 22816 12956 22880
rect 13020 22816 13036 22880
rect 13100 22816 13108 22880
rect 12788 21792 13108 22816
rect 12788 21728 12796 21792
rect 12860 21728 12876 21792
rect 12940 21728 12956 21792
rect 13020 21728 13036 21792
rect 13100 21728 13108 21792
rect 12788 20704 13108 21728
rect 12788 20640 12796 20704
rect 12860 20640 12876 20704
rect 12940 20640 12956 20704
rect 13020 20640 13036 20704
rect 13100 20640 13108 20704
rect 12788 19616 13108 20640
rect 12788 19552 12796 19616
rect 12860 19552 12876 19616
rect 12940 19552 12956 19616
rect 13020 19552 13036 19616
rect 13100 19552 13108 19616
rect 12788 18528 13108 19552
rect 12788 18464 12796 18528
rect 12860 18464 12876 18528
rect 12940 18464 12956 18528
rect 13020 18464 13036 18528
rect 13100 18464 13108 18528
rect 12788 17440 13108 18464
rect 12788 17376 12796 17440
rect 12860 17376 12876 17440
rect 12940 17376 12956 17440
rect 13020 17376 13036 17440
rect 13100 17376 13108 17440
rect 12788 16352 13108 17376
rect 12788 16288 12796 16352
rect 12860 16288 12876 16352
rect 12940 16288 12956 16352
rect 13020 16288 13036 16352
rect 13100 16288 13108 16352
rect 12788 15264 13108 16288
rect 12788 15200 12796 15264
rect 12860 15200 12876 15264
rect 12940 15200 12956 15264
rect 13020 15200 13036 15264
rect 13100 15200 13108 15264
rect 12788 14176 13108 15200
rect 12788 14112 12796 14176
rect 12860 14112 12876 14176
rect 12940 14112 12956 14176
rect 13020 14112 13036 14176
rect 13100 14112 13108 14176
rect 12788 13088 13108 14112
rect 12788 13024 12796 13088
rect 12860 13024 12876 13088
rect 12940 13024 12956 13088
rect 13020 13024 13036 13088
rect 13100 13024 13108 13088
rect 12788 12000 13108 13024
rect 12788 11936 12796 12000
rect 12860 11936 12876 12000
rect 12940 11936 12956 12000
rect 13020 11936 13036 12000
rect 13100 11936 13108 12000
rect 12788 10912 13108 11936
rect 12788 10848 12796 10912
rect 12860 10848 12876 10912
rect 12940 10848 12956 10912
rect 13020 10848 13036 10912
rect 13100 10848 13108 10912
rect 12788 9824 13108 10848
rect 12788 9760 12796 9824
rect 12860 9760 12876 9824
rect 12940 9760 12956 9824
rect 13020 9760 13036 9824
rect 13100 9760 13108 9824
rect 12788 8736 13108 9760
rect 12788 8672 12796 8736
rect 12860 8672 12876 8736
rect 12940 8672 12956 8736
rect 13020 8672 13036 8736
rect 13100 8672 13108 8736
rect 11283 8396 11349 8397
rect 11283 8332 11284 8396
rect 11348 8332 11349 8396
rect 11283 8331 11349 8332
rect 10814 8128 10822 8192
rect 10886 8128 10902 8192
rect 10966 8128 10982 8192
rect 11046 8128 11062 8192
rect 11126 8128 11134 8192
rect 10547 8124 10613 8125
rect 10547 8060 10548 8124
rect 10612 8060 10613 8124
rect 10547 8059 10613 8060
rect 10363 7852 10429 7853
rect 10363 7788 10364 7852
rect 10428 7788 10429 7852
rect 10363 7787 10429 7788
rect 10179 7716 10245 7717
rect 10179 7652 10180 7716
rect 10244 7652 10245 7716
rect 10179 7651 10245 7652
rect 9995 7580 10061 7581
rect 9995 7516 9996 7580
rect 10060 7516 10061 7580
rect 9995 7515 10061 7516
rect 10814 7104 11134 8128
rect 10814 7040 10822 7104
rect 10886 7040 10902 7104
rect 10966 7040 10982 7104
rect 11046 7040 11062 7104
rect 11126 7040 11134 7104
rect 10814 6016 11134 7040
rect 10814 5952 10822 6016
rect 10886 5952 10902 6016
rect 10966 5952 10982 6016
rect 11046 5952 11062 6016
rect 11126 5952 11134 6016
rect 10814 4928 11134 5952
rect 11286 5133 11346 8331
rect 12788 7648 13108 8672
rect 12788 7584 12796 7648
rect 12860 7584 12876 7648
rect 12940 7584 12956 7648
rect 13020 7584 13036 7648
rect 13100 7584 13108 7648
rect 12788 6560 13108 7584
rect 12788 6496 12796 6560
rect 12860 6496 12876 6560
rect 12940 6496 12956 6560
rect 13020 6496 13036 6560
rect 13100 6496 13108 6560
rect 12788 5472 13108 6496
rect 12788 5408 12796 5472
rect 12860 5408 12876 5472
rect 12940 5408 12956 5472
rect 13020 5408 13036 5472
rect 13100 5408 13108 5472
rect 11283 5132 11349 5133
rect 11283 5068 11284 5132
rect 11348 5068 11349 5132
rect 11283 5067 11349 5068
rect 10814 4864 10822 4928
rect 10886 4864 10902 4928
rect 10966 4864 10982 4928
rect 11046 4864 11062 4928
rect 11126 4864 11134 4928
rect 10814 3840 11134 4864
rect 10814 3776 10822 3840
rect 10886 3776 10902 3840
rect 10966 3776 10982 3840
rect 11046 3776 11062 3840
rect 11126 3776 11134 3840
rect 9811 3092 9877 3093
rect 9811 3028 9812 3092
rect 9876 3028 9877 3092
rect 9811 3027 9877 3028
rect 8840 2144 8848 2208
rect 8912 2144 8928 2208
rect 8992 2144 9008 2208
rect 9072 2144 9088 2208
rect 9152 2144 9160 2208
rect 8840 1120 9160 2144
rect 8840 1056 8848 1120
rect 8912 1056 8928 1120
rect 8992 1056 9008 1120
rect 9072 1056 9088 1120
rect 9152 1056 9160 1120
rect 8840 1040 9160 1056
rect 10814 2752 11134 3776
rect 10814 2688 10822 2752
rect 10886 2688 10902 2752
rect 10966 2688 10982 2752
rect 11046 2688 11062 2752
rect 11126 2688 11134 2752
rect 10814 1664 11134 2688
rect 10814 1600 10822 1664
rect 10886 1600 10902 1664
rect 10966 1600 10982 1664
rect 11046 1600 11062 1664
rect 11126 1600 11134 1664
rect 10814 1040 11134 1600
rect 12788 4384 13108 5408
rect 12788 4320 12796 4384
rect 12860 4320 12876 4384
rect 12940 4320 12956 4384
rect 13020 4320 13036 4384
rect 13100 4320 13108 4384
rect 12788 3296 13108 4320
rect 12788 3232 12796 3296
rect 12860 3232 12876 3296
rect 12940 3232 12956 3296
rect 13020 3232 13036 3296
rect 13100 3232 13108 3296
rect 12788 2208 13108 3232
rect 12788 2144 12796 2208
rect 12860 2144 12876 2208
rect 12940 2144 12956 2208
rect 13020 2144 13036 2208
rect 13100 2144 13108 2208
rect 12788 1120 13108 2144
rect 12788 1056 12796 1120
rect 12860 1056 12876 1120
rect 12940 1056 12956 1120
rect 13020 1056 13036 1120
rect 13100 1056 13108 1120
rect 12788 1040 13108 1056
rect 14762 22336 15082 22896
rect 14762 22272 14770 22336
rect 14834 22272 14850 22336
rect 14914 22272 14930 22336
rect 14994 22272 15010 22336
rect 15074 22272 15082 22336
rect 14762 21248 15082 22272
rect 14762 21184 14770 21248
rect 14834 21184 14850 21248
rect 14914 21184 14930 21248
rect 14994 21184 15010 21248
rect 15074 21184 15082 21248
rect 14762 20160 15082 21184
rect 14762 20096 14770 20160
rect 14834 20096 14850 20160
rect 14914 20096 14930 20160
rect 14994 20096 15010 20160
rect 15074 20096 15082 20160
rect 14762 19072 15082 20096
rect 14762 19008 14770 19072
rect 14834 19008 14850 19072
rect 14914 19008 14930 19072
rect 14994 19008 15010 19072
rect 15074 19008 15082 19072
rect 14762 17984 15082 19008
rect 14762 17920 14770 17984
rect 14834 17920 14850 17984
rect 14914 17920 14930 17984
rect 14994 17920 15010 17984
rect 15074 17920 15082 17984
rect 14762 16896 15082 17920
rect 14762 16832 14770 16896
rect 14834 16832 14850 16896
rect 14914 16832 14930 16896
rect 14994 16832 15010 16896
rect 15074 16832 15082 16896
rect 14762 15808 15082 16832
rect 14762 15744 14770 15808
rect 14834 15744 14850 15808
rect 14914 15744 14930 15808
rect 14994 15744 15010 15808
rect 15074 15744 15082 15808
rect 14762 14720 15082 15744
rect 14762 14656 14770 14720
rect 14834 14656 14850 14720
rect 14914 14656 14930 14720
rect 14994 14656 15010 14720
rect 15074 14656 15082 14720
rect 14762 13632 15082 14656
rect 14762 13568 14770 13632
rect 14834 13568 14850 13632
rect 14914 13568 14930 13632
rect 14994 13568 15010 13632
rect 15074 13568 15082 13632
rect 14762 12544 15082 13568
rect 14762 12480 14770 12544
rect 14834 12480 14850 12544
rect 14914 12480 14930 12544
rect 14994 12480 15010 12544
rect 15074 12480 15082 12544
rect 14762 11456 15082 12480
rect 14762 11392 14770 11456
rect 14834 11392 14850 11456
rect 14914 11392 14930 11456
rect 14994 11392 15010 11456
rect 15074 11392 15082 11456
rect 14762 10368 15082 11392
rect 14762 10304 14770 10368
rect 14834 10304 14850 10368
rect 14914 10304 14930 10368
rect 14994 10304 15010 10368
rect 15074 10304 15082 10368
rect 14762 9280 15082 10304
rect 14762 9216 14770 9280
rect 14834 9216 14850 9280
rect 14914 9216 14930 9280
rect 14994 9216 15010 9280
rect 15074 9216 15082 9280
rect 14762 8192 15082 9216
rect 14762 8128 14770 8192
rect 14834 8128 14850 8192
rect 14914 8128 14930 8192
rect 14994 8128 15010 8192
rect 15074 8128 15082 8192
rect 14762 7104 15082 8128
rect 14762 7040 14770 7104
rect 14834 7040 14850 7104
rect 14914 7040 14930 7104
rect 14994 7040 15010 7104
rect 15074 7040 15082 7104
rect 14762 6016 15082 7040
rect 14762 5952 14770 6016
rect 14834 5952 14850 6016
rect 14914 5952 14930 6016
rect 14994 5952 15010 6016
rect 15074 5952 15082 6016
rect 14762 4928 15082 5952
rect 14762 4864 14770 4928
rect 14834 4864 14850 4928
rect 14914 4864 14930 4928
rect 14994 4864 15010 4928
rect 15074 4864 15082 4928
rect 14762 3840 15082 4864
rect 14762 3776 14770 3840
rect 14834 3776 14850 3840
rect 14914 3776 14930 3840
rect 14994 3776 15010 3840
rect 15074 3776 15082 3840
rect 14762 2752 15082 3776
rect 14762 2688 14770 2752
rect 14834 2688 14850 2752
rect 14914 2688 14930 2752
rect 14994 2688 15010 2752
rect 15074 2688 15082 2752
rect 14762 1664 15082 2688
rect 14762 1600 14770 1664
rect 14834 1600 14850 1664
rect 14914 1600 14930 1664
rect 14994 1600 15010 1664
rect 15074 1600 15082 1664
rect 14762 1040 15082 1600
use sky130_ef_sc_hd__decap_12  FILLER_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_25
timestamp 1649977179
transform 1 0 3404 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_37
timestamp 1649977179
transform 1 0 4508 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5612 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1649977179
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1649977179
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1649977179
transform 1 0 2116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_22
timestamp 1649977179
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_29
timestamp 1649977179
transform 1 0 3772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_41
timestamp 1649977179
transform 1 0 4876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_16
timestamp 1649977179
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1649977179
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1649977179
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_39
timestamp 1649977179
transform 1 0 4692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_51
timestamp 1649977179
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_63
timestamp 1649977179
transform 1 0 6900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1649977179
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1649977179
transform 1 0 3220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1649977179
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_46
timestamp 1649977179
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_35
timestamp 1649977179
transform 1 0 4324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_49
timestamp 1649977179
transform 1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_56
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_63
timestamp 1649977179
transform 1 0 6900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1649977179
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1649977179
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_28
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1649977179
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_67
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_79
timestamp 1649977179
transform 1 0 8372 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_91
timestamp 1649977179
transform 1 0 9476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp 1649977179
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_18
timestamp 1649977179
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_39
timestamp 1649977179
transform 1 0 4692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_50
timestamp 1649977179
transform 1 0 5704 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_59
timestamp 1649977179
transform 1 0 6532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_66
timestamp 1649977179
transform 1 0 7176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_73
timestamp 1649977179
transform 1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 1649977179
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_33
timestamp 1649977179
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_44
timestamp 1649977179
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_63
timestamp 1649977179
transform 1 0 6900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_72
timestamp 1649977179
transform 1 0 7728 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_79
timestamp 1649977179
transform 1 0 8372 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_86
timestamp 1649977179
transform 1 0 9016 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_98
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_39
timestamp 1649977179
transform 1 0 4692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_50
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_61
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_71
timestamp 1649977179
transform 1 0 7636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1649977179
transform 1 0 9200 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_95
timestamp 1649977179
transform 1 0 9844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_107
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_119
timestamp 1649977179
transform 1 0 12052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1649977179
transform 1 0 13156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1649977179
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_44
timestamp 1649977179
transform 1 0 5152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_64
timestamp 1649977179
transform 1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_75
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_98
timestamp 1649977179
transform 1 0 10120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1649977179
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_49
timestamp 1649977179
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1649977179
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_73
timestamp 1649977179
transform 1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_91
timestamp 1649977179
transform 1 0 9476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_98
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_105
timestamp 1649977179
transform 1 0 10764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_112
timestamp 1649977179
transform 1 0 11408 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_119
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_131
timestamp 1649977179
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_24
timestamp 1649977179
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1649977179
transform 1 0 8280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_89
timestamp 1649977179
transform 1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_116
timestamp 1649977179
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_123
timestamp 1649977179
transform 1 0 12420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_135
timestamp 1649977179
transform 1 0 13524 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_147
timestamp 1649977179
transform 1 0 14628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_159
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_49
timestamp 1649977179
transform 1 0 5612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_63
timestamp 1649977179
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_76
timestamp 1649977179
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_92
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_103
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_112
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_119
timestamp 1649977179
transform 1 0 12052 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_126
timestamp 1649977179
transform 1 0 12696 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_25
timestamp 1649977179
transform 1 0 3404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1649977179
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_73
timestamp 1649977179
transform 1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_85
timestamp 1649977179
transform 1 0 8924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_97
timestamp 1649977179
transform 1 0 10028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1649977179
transform 1 0 11960 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_126
timestamp 1649977179
transform 1 0 12696 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_133
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1649977179
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_78
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_94
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_106
timestamp 1649977179
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_127
timestamp 1649977179
transform 1 0 12788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_134
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_144
timestamp 1649977179
transform 1 0 14352 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_156
timestamp 1649977179
transform 1 0 15456 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_23
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_104
timestamp 1649977179
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_119
timestamp 1649977179
transform 1 0 12052 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1649977179
transform 1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_134
timestamp 1649977179
transform 1 0 13432 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_141
timestamp 1649977179
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_148
timestamp 1649977179
transform 1 0 14720 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1649977179
transform 1 0 8280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_94
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_122
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_129
timestamp 1649977179
transform 1 0 12972 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1649977179
transform 1 0 3772 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1649977179
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_73
timestamp 1649977179
transform 1 0 7820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_85
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_116
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_123
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_135
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_147
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_50
timestamp 1649977179
transform 1 0 5704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_70
timestamp 1649977179
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_91
timestamp 1649977179
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1649977179
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1649977179
transform 1 0 11592 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_6
timestamp 1649977179
transform 1 0 1656 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_31
timestamp 1649977179
transform 1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_73
timestamp 1649977179
transform 1 0 7820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_83
timestamp 1649977179
transform 1 0 8740 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_92
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1649977179
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1649977179
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1649977179
transform 1 0 5244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1649977179
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_89
timestamp 1649977179
transform 1 0 9292 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_96
timestamp 1649977179
transform 1 0 9936 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_108
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_120
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_132
timestamp 1649977179
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_23
timestamp 1649977179
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1649977179
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_66
timestamp 1649977179
transform 1 0 7176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_76
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_83
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_90
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_102
timestamp 1649977179
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_58
timestamp 1649977179
transform 1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 1649977179
transform 1 0 7544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_23
timestamp 1649977179
transform 1 0 3220 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1649977179
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_61
timestamp 1649977179
transform 1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_68
timestamp 1649977179
transform 1 0 7360 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_80
timestamp 1649977179
transform 1 0 8464 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_92
timestamp 1649977179
transform 1 0 9568 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_104
timestamp 1649977179
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1649977179
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_39
timestamp 1649977179
transform 1 0 4692 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_50
timestamp 1649977179
transform 1 0 5704 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_57
timestamp 1649977179
transform 1 0 6348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_69
timestamp 1649977179
transform 1 0 7452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1649977179
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_19
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1649977179
transform 1 0 4140 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1649977179
transform 1 0 5244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1649977179
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1649977179
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_33
timestamp 1649977179
transform 1 0 4140 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_40
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_52
timestamp 1649977179
transform 1 0 5888 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_64
timestamp 1649977179
transform 1 0 6992 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_76
timestamp 1649977179
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_16
timestamp 1649977179
transform 1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_24
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1649977179
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1649977179
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_14
timestamp 1649977179
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_26
timestamp 1649977179
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_38
timestamp 1649977179
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_50
timestamp 1649977179
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_14
timestamp 1649977179
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1649977179
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_7
timestamp 1649977179
transform 1 0 1748 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_19
timestamp 1649977179
transform 1 0 2852 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_31
timestamp 1649977179
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1649977179
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_29
timestamp 1649977179
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_41
timestamp 1649977179
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1649977179
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_85
timestamp 1649977179
transform 1 0 8924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_97
timestamp 1649977179
transform 1 0 10028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1649977179
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_141
timestamp 1649977179
transform 1 0 14076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_153
timestamp 1649977179
transform 1 0 15180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1649977179
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 16836 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 16836 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 16836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 16836 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 16836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 16836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 16836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 16836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 3680 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 8832 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 13984 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9936 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4692 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _118_
timestamp 1649977179
transform -1 0 4140 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _119_
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14076 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1649977179
transform -1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _123_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9292 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8464 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9568 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1649977179
transform -1 0 7360 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _128_
timestamp 1649977179
transform 1 0 5336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1649977179
transform 1 0 11776 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1649977179
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _131_
timestamp 1649977179
transform 1 0 12144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1649977179
transform -1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _134_
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 1649977179
transform -1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8740 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp 1649977179
transform -1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _140_
timestamp 1649977179
transform 1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _141_
timestamp 1649977179
transform 1 0 5060 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7452 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _143_
timestamp 1649977179
transform -1 0 4140 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _144_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5704 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _145_
timestamp 1649977179
transform 1 0 11316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1649977179
transform 1 0 12696 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _147_
timestamp 1649977179
transform -1 0 3772 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1649977179
transform 1 0 12052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _150_
timestamp 1649977179
transform -1 0 3312 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1649977179
transform 1 0 8464 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _153_
timestamp 1649977179
transform -1 0 3956 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _155_
timestamp 1649977179
transform -1 0 12236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7452 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _158_
timestamp 1649977179
transform -1 0 2484 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _160_
timestamp 1649977179
transform 1 0 5612 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _161_
timestamp 1649977179
transform -1 0 8464 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6808 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5060 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _165_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp 1649977179
transform -1 0 2576 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1649977179
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _168_
timestamp 1649977179
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _170_
timestamp 1649977179
transform 1 0 13064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _171_
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5888 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11868 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _174_
timestamp 1649977179
transform -1 0 10120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9476 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4048 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _178_
timestamp 1649977179
transform 1 0 5060 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7268 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _180_
timestamp 1649977179
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _181_
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _183_
timestamp 1649977179
transform -1 0 9752 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _184_
timestamp 1649977179
transform -1 0 9476 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10212 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _186_
timestamp 1649977179
transform 1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _187_
timestamp 1649977179
transform -1 0 4324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _188_
timestamp 1649977179
transform -1 0 8924 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _189_
timestamp 1649977179
transform -1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _190_
timestamp 1649977179
transform 1 0 2668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10764 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _192_
timestamp 1649977179
transform 1 0 5428 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _193_
timestamp 1649977179
transform 1 0 8188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _194_
timestamp 1649977179
transform -1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1649977179
transform 1 0 13156 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _196_
timestamp 1649977179
transform 1 0 5520 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _197_
timestamp 1649977179
transform -1 0 11960 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _198_
timestamp 1649977179
transform -1 0 7636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10856 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _200_
timestamp 1649977179
transform 1 0 10028 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _201_
timestamp 1649977179
transform -1 0 11684 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12788 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _203_
timestamp 1649977179
transform 1 0 4508 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _204_
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _205_
timestamp 1649977179
transform 1 0 10396 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9292 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _208_
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _209_
timestamp 1649977179
transform 1 0 2852 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _210_
timestamp 1649977179
transform -1 0 9568 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _211_
timestamp 1649977179
transform 1 0 7544 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _212_
timestamp 1649977179
transform 1 0 10948 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _213_
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _214_
timestamp 1649977179
transform 1 0 7544 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _216_
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _217_
timestamp 1649977179
transform -1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _218_
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _219_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _220_
timestamp 1649977179
transform 1 0 9292 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9476 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1649977179
transform 1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _223_
timestamp 1649977179
transform 1 0 2668 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _224_
timestamp 1649977179
transform 1 0 6072 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _227_
timestamp 1649977179
transform -1 0 5520 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _229_
timestamp 1649977179
transform -1 0 7728 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 1649977179
transform 1 0 5612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _231_
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _232_
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _233_
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1649977179
transform -1 0 7176 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _235_
timestamp 1649977179
transform 1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1649977179
transform -1 0 6808 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _238_
timestamp 1649977179
transform -1 0 9752 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp 1649977179
transform 1 0 9660 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _240_
timestamp 1649977179
transform -1 0 10580 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _241_
timestamp 1649977179
transform -1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _242_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _244_
timestamp 1649977179
transform -1 0 2668 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _245_
timestamp 1649977179
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _246_
timestamp 1649977179
transform -1 0 10120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _247_
timestamp 1649977179
transform -1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _248_
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _249_
timestamp 1649977179
transform -1 0 12420 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _250_
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _251_
timestamp 1649977179
transform -1 0 2760 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _252_
timestamp 1649977179
transform -1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _253_
timestamp 1649977179
transform -1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp 1649977179
transform -1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _255_
timestamp 1649977179
transform -1 0 12696 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _256_
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _257_
timestamp 1649977179
transform -1 0 12052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp 1649977179
transform 1 0 2024 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _259_
timestamp 1649977179
transform -1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1472 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _261_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _262_
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _263_
timestamp 1649977179
transform 1 0 1472 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _265_
timestamp 1649977179
transform 1 0 3680 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _266_
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _267_
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _268_
timestamp 1649977179
transform -1 0 3312 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _269_
timestamp 1649977179
transform -1 0 3312 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _270_
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _271_
timestamp 1649977179
transform -1 0 5612 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3404 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _274_
timestamp 1649977179
transform -1 0 5244 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _275_
timestamp 1649977179
transform -1 0 7084 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _276_
timestamp 1649977179
transform -1 0 5244 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _277_
timestamp 1649977179
transform -1 0 7084 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _278_
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _279_
timestamp 1649977179
transform 1 0 1656 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _280_
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _281_
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _282_
timestamp 1649977179
transform -1 0 5612 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _283_
timestamp 1649977179
transform -1 0 5244 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _284_
timestamp 1649977179
transform -1 0 5060 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _285_
timestamp 1649977179
transform -1 0 7544 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _286_
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _287_
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _288_
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _289_
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _290_
timestamp 1649977179
transform -1 0 7820 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _291_
timestamp 1649977179
transform -1 0 2852 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _292_
timestamp 1649977179
transform -1 0 7820 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _293_
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _294_
timestamp 1649977179
transform 1 0 3680 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _295_
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _296_
timestamp 1649977179
transform 1 0 5612 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _297_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _298_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _300_
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _301_
timestamp 1649977179
transform -1 0 4140 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _302_
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _303_
timestamp 1649977179
transform 1 0 2116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _304_
timestamp 1649977179
transform -1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _305_
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _306_
timestamp 1649977179
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 1656 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 1656 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater7
timestamp 1649977179
transform -1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater8
timestamp 1649977179
transform 1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater9
timestamp 1649977179
transform -1 0 2944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater10
timestamp 1649977179
transform -1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater11
timestamp 1649977179
transform -1 0 6900 0 1 4352
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 688 400 808 0 FreeSans 480 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 0 2184 400 2304 0 FreeSans 480 0 0 0 io_in[1]
port 1 nsew signal input
flabel metal3 s 0 3680 400 3800 0 FreeSans 480 0 0 0 io_in[2]
port 2 nsew signal input
flabel metal3 s 0 5176 400 5296 0 FreeSans 480 0 0 0 io_in[3]
port 3 nsew signal input
flabel metal3 s 0 6672 400 6792 0 FreeSans 480 0 0 0 io_in[4]
port 4 nsew signal input
flabel metal3 s 0 8168 400 8288 0 FreeSans 480 0 0 0 io_in[5]
port 5 nsew signal input
flabel metal3 s 0 9664 400 9784 0 FreeSans 480 0 0 0 io_in[6]
port 6 nsew signal input
flabel metal3 s 0 11160 400 11280 0 FreeSans 480 0 0 0 io_in[7]
port 7 nsew signal input
flabel metal3 s 0 12656 400 12776 0 FreeSans 480 0 0 0 io_out[0]
port 8 nsew signal tristate
flabel metal3 s 0 14152 400 14272 0 FreeSans 480 0 0 0 io_out[1]
port 9 nsew signal tristate
flabel metal3 s 0 15648 400 15768 0 FreeSans 480 0 0 0 io_out[2]
port 10 nsew signal tristate
flabel metal3 s 0 17144 400 17264 0 FreeSans 480 0 0 0 io_out[3]
port 11 nsew signal tristate
flabel metal3 s 0 18640 400 18760 0 FreeSans 480 0 0 0 io_out[4]
port 12 nsew signal tristate
flabel metal3 s 0 20136 400 20256 0 FreeSans 480 0 0 0 io_out[5]
port 13 nsew signal tristate
flabel metal3 s 0 21632 400 21752 0 FreeSans 480 0 0 0 io_out[6]
port 14 nsew signal tristate
flabel metal3 s 0 23128 400 23248 0 FreeSans 480 0 0 0 io_out[7]
port 15 nsew signal tristate
flabel metal4 s 2918 1040 3238 22896 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 6866 1040 7186 22896 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 10814 1040 11134 22896 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 14762 1040 15082 22896 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 4892 1040 5212 22896 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 8840 1040 9160 22896 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 12788 1040 13108 22896 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 18000 24000
<< end >>
