module tholin_avalonsemi_5401 (vccd1,
    vssd1,
    io_in,
    io_out);
 input vccd1;
 input vssd1;
 input [7:0] io_in;
 output [7:0] io_out;

 wire \CIRCUIT_0.GATES_10.input1 ;
 wire \CIRCUIT_0.GATES_10.result ;
 wire \CIRCUIT_0.GATES_11.result ;
 wire \CIRCUIT_0.GATES_28.result ;
 wire \CIRCUIT_0.GATES_29.result ;
 wire \CIRCUIT_0.GATES_31.result ;
 wire \CIRCUIT_0.GATES_36.result ;
 wire \CIRCUIT_0.GATES_39.result ;
 wire \CIRCUIT_0.GATES_40.result ;
 wire \CIRCUIT_0.GATES_41.result ;
 wire \CIRCUIT_0.GATES_42.result ;
 wire \CIRCUIT_0.GATES_43.result ;
 wire \CIRCUIT_0.GATES_59.result ;
 wire \CIRCUIT_0.GATES_65.result ;
 wire \CIRCUIT_0.GATES_72.result ;
 wire \CIRCUIT_0.MEMORY_100.s_currentState ;
 wire \CIRCUIT_0.MEMORY_74.d ;
 wire \CIRCUIT_0.MEMORY_74.s_currentState ;
 wire \CIRCUIT_0.MEMORY_75.d ;
 wire \CIRCUIT_0.MEMORY_75.s_currentState ;
 wire \CIRCUIT_0.MEMORY_76.d ;
 wire \CIRCUIT_0.MEMORY_76.s_currentState ;
 wire \CIRCUIT_0.MEMORY_77.d ;
 wire \CIRCUIT_0.MEMORY_77.s_currentState ;
 wire \CIRCUIT_0.MEMORY_78.d ;
 wire \CIRCUIT_0.MEMORY_78.s_currentState ;
 wire \CIRCUIT_0.MEMORY_79.d ;
 wire \CIRCUIT_0.MEMORY_79.s_currentState ;
 wire \CIRCUIT_0.MEMORY_80.s_currentState ;
 wire \CIRCUIT_0.MEMORY_81.s_currentState ;
 wire \CIRCUIT_0.MEMORY_82.s_currentState ;
 wire \CIRCUIT_0.MEMORY_83.s_currentState ;
 wire \CIRCUIT_0.MEMORY_84.s_currentState ;
 wire \CIRCUIT_0.MEMORY_85.s_currentState ;
 wire \CIRCUIT_0.MEMORY_86.s_currentState ;
 wire \CIRCUIT_0.MEMORY_87.s_currentState ;
 wire \CIRCUIT_0.MEMORY_88.s_currentState ;
 wire \CIRCUIT_0.MEMORY_89.s_currentState ;
 wire \CIRCUIT_0.MEMORY_90.s_currentState ;
 wire \CIRCUIT_0.MEMORY_91.s_currentState ;
 wire \CIRCUIT_0.MEMORY_92.s_currentState ;
 wire \CIRCUIT_0.MEMORY_93.s_currentState ;
 wire \CIRCUIT_0.MEMORY_94.s_currentState ;
 wire \CIRCUIT_0.MEMORY_95.s_currentState ;
 wire \CIRCUIT_0.MEMORY_96.s_currentState ;
 wire \CIRCUIT_0.MEMORY_97.s_currentState ;
 wire \CIRCUIT_0.MEMORY_98.s_currentState ;
 wire \CIRCUIT_0.MEMORY_99.s_currentState ;
 wire \CIRCUIT_0.O_4_MAR ;
 wire \CIRCUIT_0.O_5_WRITE ;
 wire \CIRCUIT_0.O_6_JMP ;
 wire \CIRCUIT_0.O_7_I ;
 wire \CIRCUIT_0.O_D0_RR0 ;
 wire \CIRCUIT_0.O_D1_RR1 ;
 wire \CIRCUIT_0.O_D2_RR2 ;
 wire \CIRCUIT_0.O_D3_RR3 ;
 wire \CIRCUIT_0.dest_reg_sel_1.CLK1 ;
 wire \CIRCUIT_0.dest_reg_sel_1.GATES_1.result ;
 wire \CIRCUIT_0.dest_reg_sel_1.MEMORY_2.s_currentState ;
 wire \CIRCUIT_0.dest_reg_sel_1.MEMORY_3.s_currentState ;
 wire \CIRCUIT_0.dest_reg_sel_1.MEMORY_4.s_currentState ;
 wire \CIRCUIT_0.inst_dec_1.MEMORY_21.s_currentState ;
 wire \CIRCUIT_0.inst_dec_1.MEMORY_22.s_currentState ;
 wire \CIRCUIT_0.inst_dec_1.MEMORY_23.s_currentState ;
 wire \CIRCUIT_0.inst_dec_1.MEMORY_24.s_currentState ;
 wire \CIRCUIT_0.multiply_1.GATES_23.input2 ;
 wire \CIRCUIT_0.multiply_1.GATES_24.result ;
 wire \CIRCUIT_0.multiply_1.MEMORY_25.d ;
 wire \CIRCUIT_0.multiply_1.MEMORY_25.s_currentState ;
 wire \CIRCUIT_0.multiply_1.MEMORY_26.d ;
 wire \CIRCUIT_0.multiply_1.MEMORY_26.s_currentState ;
 wire \CIRCUIT_0.multiply_1.MEMORY_27.d ;
 wire \CIRCUIT_0.multiply_1.MEMORY_27.s_currentState ;
 wire \CIRCUIT_0.multiply_1.MEMORY_28.d ;
 wire \CIRCUIT_0.multiply_1.MEMORY_28.s_currentState ;
 wire \CIRCUIT_0.multiply_1.MEMORY_29.d ;
 wire \CIRCUIT_0.multiply_1.MEMORY_29.s_currentState ;
 wire \CIRCUIT_0.multiply_1.MEMORY_30.d ;
 wire \CIRCUIT_0.multiply_1.MEMORY_30.s_currentState ;
 wire \CIRCUIT_0.multiply_1.MEMORY_31.d ;
 wire \CIRCUIT_0.multiply_1.MEMORY_31.s_currentState ;
 wire \CIRCUIT_0.multiply_1.MEMORY_32.d ;
 wire \CIRCUIT_0.multiply_1.MEMORY_32.s_currentState ;
 wire \CIRCUIT_0.multiply_1.MEMORY_33.d ;
 wire \CIRCUIT_0.multiply_1.MEMORY_33.s_currentState ;
 wire \CIRCUIT_0.multiply_1.MEMORY_34.d ;
 wire \CIRCUIT_0.multiply_1.MEMORY_34.s_currentState ;
 wire \CIRCUIT_0.multiply_1.MEMORY_35.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_10.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_11.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_12.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_9.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_10.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_11.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_12.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_13.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_14.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_15.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_16.s_currentState ;
 wire \CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_9.s_currentState ;
 wire \CIRCUIT_0.output_logic_1.GATES_13.input2 ;
 wire \CIRCUIT_0.toggle_1.GATES_10.input1 ;
 wire \CIRCUIT_0.toggle_1.GATES_10.input2 ;
 wire \CIRCUIT_0.toggle_1.GATES_12.input1 ;
 wire \CIRCUIT_0.toggle_1.GATES_8.result ;
 wire \CIRCUIT_0.toggle_1.MEMORY_17.s_currentState ;
 wire \CIRCUIT_0.toggle_1.MEMORY_18.s_currentState ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire clknet_0__009_;
 wire clknet_0__218_;
 wire clknet_0__226_;
 wire clknet_0__227_;
 wire clknet_1_0__leaf__009_;
 wire clknet_1_0__leaf__218_;
 wire clknet_1_0__leaf__226_;
 wire clknet_1_0__leaf__227_;
 wire clknet_1_1__leaf__009_;
 wire clknet_1_1__leaf__218_;
 wire clknet_1_1__leaf__226_;
 wire clknet_1_1__leaf__227_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire [0:0] clknet_0_io_in;
 wire [0:0] clknet_1_0__leaf_io_in;
 wire [0:0] clknet_1_1__leaf_io_in;

 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 _238_ (.A(\CIRCUIT_0.MEMORY_80.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_047_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(\CIRCUIT_0.GATES_59.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_000_));
 sky130_fd_sc_hd__or2_1 _240_ (.A(_047_),
    .B(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_048_));
 sky130_fd_sc_hd__clkbuf_1 _241_ (.A(\CIRCUIT_0.MEMORY_75.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_049_));
 sky130_fd_sc_hd__and3b_1 _242_ (.A_N(\CIRCUIT_0.inst_dec_1.MEMORY_22.s_currentState ),
    .B(\CIRCUIT_0.MEMORY_86.s_currentState ),
    .C(\CIRCUIT_0.MEMORY_87.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_050_));
 sky130_fd_sc_hd__and4bb_1 _243_ (.A_N(\CIRCUIT_0.inst_dec_1.MEMORY_24.s_currentState ),
    .B_N(\CIRCUIT_0.inst_dec_1.MEMORY_23.s_currentState ),
    .C(\CIRCUIT_0.MEMORY_85.s_currentState ),
    .D(\CIRCUIT_0.MEMORY_84.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_051_));
 sky130_fd_sc_hd__nand3_1 _244_ (.A(\CIRCUIT_0.MEMORY_81.s_currentState ),
    .B(_050_),
    .C(_051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_052_));
 sky130_fd_sc_hd__nor2_1 _245_ (.A(\CIRCUIT_0.MEMORY_83.s_currentState ),
    .B(\CIRCUIT_0.MEMORY_82.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_053_));
 sky130_fd_sc_hd__and4_1 _246_ (.A(\CIRCUIT_0.MEMORY_81.s_currentState ),
    .B(_050_),
    .C(_051_),
    .D(_053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _247_ (.A0(\CIRCUIT_0.multiply_1.MEMORY_32.s_currentState ),
    .A1(\CIRCUIT_0.multiply_1.MEMORY_28.s_currentState ),
    .S(_047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_055_));
 sky130_fd_sc_hd__a22o_1 _248_ (.A1(net5),
    .A2(_052_),
    .B1(_054_),
    .B2(_055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _249_ (.A0(_049_),
    .A1(_056_),
    .S(\CIRCUIT_0.MEMORY_74.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_057_));
 sky130_fd_sc_hd__clkbuf_1 _250_ (.A(_057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.GATES_36.result ));
 sky130_fd_sc_hd__or2_1 _251_ (.A(_048_),
    .B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_058_));
 sky130_fd_sc_hd__clkbuf_1 _252_ (.A(_058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_036_));
 sky130_fd_sc_hd__clkbuf_1 _253_ (.A(\CIRCUIT_0.MEMORY_79.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _254_ (.A0(\CIRCUIT_0.multiply_1.MEMORY_31.s_currentState ),
    .A1(\CIRCUIT_0.multiply_1.MEMORY_27.s_currentState ),
    .S(\CIRCUIT_0.MEMORY_80.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_060_));
 sky130_fd_sc_hd__a22o_1 _255_ (.A1(net4),
    .A2(_052_),
    .B1(_054_),
    .B2(_060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _256_ (.A0(_059_),
    .A1(_061_),
    .S(\CIRCUIT_0.MEMORY_74.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_062_));
 sky130_fd_sc_hd__clkbuf_1 _257_ (.A(_062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.GATES_31.result ));
 sky130_fd_sc_hd__or2_1 _258_ (.A(_048_),
    .B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_063_));
 sky130_fd_sc_hd__clkbuf_1 _259_ (.A(_063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_034_));
 sky130_fd_sc_hd__clkbuf_1 _260_ (.A(\CIRCUIT_0.MEMORY_78.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _261_ (.A0(\CIRCUIT_0.multiply_1.MEMORY_30.s_currentState ),
    .A1(\CIRCUIT_0.multiply_1.MEMORY_26.s_currentState ),
    .S(\CIRCUIT_0.MEMORY_80.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_065_));
 sky130_fd_sc_hd__and4_1 _262_ (.A(\CIRCUIT_0.MEMORY_80.s_currentState ),
    .B(\CIRCUIT_0.MEMORY_81.s_currentState ),
    .C(\CIRCUIT_0.MEMORY_83.s_currentState ),
    .D(\CIRCUIT_0.MEMORY_82.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_066_));
 sky130_fd_sc_hd__and4_1 _263_ (.A(net7),
    .B(_050_),
    .C(_051_),
    .D(_066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_067_));
 sky130_fd_sc_hd__a221o_1 _264_ (.A1(net3),
    .A2(_052_),
    .B1(_054_),
    .B2(_065_),
    .C1(_067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _265_ (.A0(_064_),
    .A1(_068_),
    .S(\CIRCUIT_0.MEMORY_74.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_069_));
 sky130_fd_sc_hd__clkbuf_1 _266_ (.A(_069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.GATES_29.result ));
 sky130_fd_sc_hd__or2_1 _267_ (.A(_048_),
    .B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_070_));
 sky130_fd_sc_hd__clkbuf_1 _268_ (.A(_070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _269_ (.A0(\CIRCUIT_0.multiply_1.MEMORY_29.s_currentState ),
    .A1(\CIRCUIT_0.multiply_1.MEMORY_25.s_currentState ),
    .S(\CIRCUIT_0.MEMORY_80.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_071_));
 sky130_fd_sc_hd__and4_1 _270_ (.A(net6),
    .B(_050_),
    .C(_051_),
    .D(_066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_072_));
 sky130_fd_sc_hd__a221o_1 _271_ (.A1(net2),
    .A2(_052_),
    .B1(_054_),
    .B2(_071_),
    .C1(_072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _272_ (.A0(\CIRCUIT_0.MEMORY_77.s_currentState ),
    .A1(_073_),
    .S(\CIRCUIT_0.MEMORY_74.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_1 _273_ (.A(_074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.GATES_28.result ));
 sky130_fd_sc_hd__or2_1 _274_ (.A(_048_),
    .B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _275_ (.A(_075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_030_));
 sky130_fd_sc_hd__and2_1 _276_ (.A(_047_),
    .B(\CIRCUIT_0.GATES_59.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_076_));
 sky130_fd_sc_hd__clkbuf_1 _277_ (.A(_076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.multiply_1.GATES_24.result ));
 sky130_fd_sc_hd__inv_2 _278_ (.A(\CIRCUIT_0.multiply_1.GATES_24.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_028_));
 sky130_fd_sc_hd__clkbuf_1 _279_ (.A(\CIRCUIT_0.multiply_1.GATES_24.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_077_));
 sky130_fd_sc_hd__clkbuf_2 _280_ (.A(_077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_078_));
 sky130_fd_sc_hd__inv_2 _281_ (.A(_078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _282_ (.A(_078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _283_ (.A(_078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_022_));
 sky130_fd_sc_hd__or2_1 _284_ (.A(_028_),
    .B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_079_));
 sky130_fd_sc_hd__clkbuf_1 _285_ (.A(_079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_020_));
 sky130_fd_sc_hd__or2_1 _286_ (.A(_028_),
    .B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_080_));
 sky130_fd_sc_hd__clkbuf_1 _287_ (.A(_080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_018_));
 sky130_fd_sc_hd__or2_1 _288_ (.A(_028_),
    .B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_081_));
 sky130_fd_sc_hd__clkbuf_1 _289_ (.A(_081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_016_));
 sky130_fd_sc_hd__or2_1 _290_ (.A(_028_),
    .B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_082_));
 sky130_fd_sc_hd__clkbuf_1 _291_ (.A(_082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_014_));
 sky130_fd_sc_hd__inv_2 _292_ (.A(_078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _293_ (.A(_078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_010_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _294_ (.A(_077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_083_));
 sky130_fd_sc_hd__inv_2 _295_ (.A(_083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_008_));
 sky130_fd_sc_hd__clkbuf_1 _296_ (.A(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_12.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_084_));
 sky130_fd_sc_hd__nand3_1 _297_ (.A(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_12.s_currentState ),
    .B(\CIRCUIT_0.multiply_1.MEMORY_26.s_currentState ),
    .C(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_14.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_085_));
 sky130_fd_sc_hd__and3_1 _298_ (.A(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_12.s_currentState ),
    .B(\CIRCUIT_0.multiply_1.MEMORY_25.s_currentState ),
    .C(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_13.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_086_));
 sky130_fd_sc_hd__a21o_1 _299_ (.A1(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_12.s_currentState ),
    .A2(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_14.s_currentState ),
    .B1(\CIRCUIT_0.multiply_1.MEMORY_26.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_087_));
 sky130_fd_sc_hd__and3_1 _300_ (.A(_085_),
    .B(_086_),
    .C(_087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_088_));
 sky130_fd_sc_hd__a31o_1 _301_ (.A1(_084_),
    .A2(\CIRCUIT_0.multiply_1.MEMORY_26.s_currentState ),
    .A3(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_14.s_currentState ),
    .B1(_088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_089_));
 sky130_fd_sc_hd__a21o_1 _302_ (.A1(_084_),
    .A2(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_15.s_currentState ),
    .B1(\CIRCUIT_0.multiply_1.MEMORY_27.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_090_));
 sky130_fd_sc_hd__and3_1 _303_ (.A(_084_),
    .B(\CIRCUIT_0.multiply_1.MEMORY_27.s_currentState ),
    .C(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_15.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_091_));
 sky130_fd_sc_hd__inv_2 _304_ (.A(_091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_092_));
 sky130_fd_sc_hd__nand2_1 _305_ (.A(_090_),
    .B(_092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_093_));
 sky130_fd_sc_hd__xnor2_1 _306_ (.A(_089_),
    .B(_093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.multiply_1.MEMORY_27.d ));
 sky130_fd_sc_hd__clkbuf_1 _307_ (.A(_084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_094_));
 sky130_fd_sc_hd__a21o_1 _308_ (.A1(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_16.s_currentState ),
    .A2(_094_),
    .B1(\CIRCUIT_0.multiply_1.MEMORY_28.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_095_));
 sky130_fd_sc_hd__and3_1 _309_ (.A(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_16.s_currentState ),
    .B(_084_),
    .C(\CIRCUIT_0.multiply_1.MEMORY_28.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_096_));
 sky130_fd_sc_hd__inv_2 _310_ (.A(_096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_097_));
 sky130_fd_sc_hd__nand2_1 _311_ (.A(_095_),
    .B(_097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_098_));
 sky130_fd_sc_hd__a21o_1 _312_ (.A1(_089_),
    .A2(_090_),
    .B1(_091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_099_));
 sky130_fd_sc_hd__xnor2_1 _313_ (.A(_098_),
    .B(_099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.multiply_1.MEMORY_28.d ));
 sky130_fd_sc_hd__a21o_1 _314_ (.A1(_094_),
    .A2(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_9.s_currentState ),
    .B1(\CIRCUIT_0.multiply_1.MEMORY_29.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_100_));
 sky130_fd_sc_hd__and3_1 _315_ (.A(_094_),
    .B(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_9.s_currentState ),
    .C(\CIRCUIT_0.multiply_1.MEMORY_29.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_101_));
 sky130_fd_sc_hd__inv_2 _316_ (.A(_101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_102_));
 sky130_fd_sc_hd__nand2_1 _317_ (.A(_100_),
    .B(_102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_103_));
 sky130_fd_sc_hd__a21o_1 _318_ (.A1(_095_),
    .A2(_099_),
    .B1(_096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_104_));
 sky130_fd_sc_hd__xnor2_1 _319_ (.A(_103_),
    .B(_104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.multiply_1.MEMORY_29.d ));
 sky130_fd_sc_hd__clkbuf_1 _320_ (.A(_094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_105_));
 sky130_fd_sc_hd__a21oi_1 _321_ (.A1(_105_),
    .A2(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_10.s_currentState ),
    .B1(\CIRCUIT_0.multiply_1.MEMORY_30.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_106_));
 sky130_fd_sc_hd__and3_1 _322_ (.A(_094_),
    .B(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_10.s_currentState ),
    .C(\CIRCUIT_0.multiply_1.MEMORY_30.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_107_));
 sky130_fd_sc_hd__nor2_1 _323_ (.A(_106_),
    .B(_107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_108_));
 sky130_fd_sc_hd__a21o_1 _324_ (.A1(_100_),
    .A2(_104_),
    .B1(_101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_109_));
 sky130_fd_sc_hd__xor2_1 _325_ (.A(_108_),
    .B(_109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.multiply_1.MEMORY_30.d ));
 sky130_fd_sc_hd__a21oi_1 _326_ (.A1(_105_),
    .A2(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_11.s_currentState ),
    .B1(\CIRCUIT_0.multiply_1.MEMORY_31.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_110_));
 sky130_fd_sc_hd__and3_1 _327_ (.A(_105_),
    .B(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_11.s_currentState ),
    .C(\CIRCUIT_0.multiply_1.MEMORY_31.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_111_));
 sky130_fd_sc_hd__nor2_1 _328_ (.A(_110_),
    .B(_111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_112_));
 sky130_fd_sc_hd__a21o_1 _329_ (.A1(_108_),
    .A2(_109_),
    .B1(_107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_113_));
 sky130_fd_sc_hd__xor2_1 _330_ (.A(_112_),
    .B(_113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.multiply_1.MEMORY_31.d ));
 sky130_fd_sc_hd__a21o_1 _331_ (.A1(_112_),
    .A2(_113_),
    .B1(_111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_114_));
 sky130_fd_sc_hd__nand2_1 _332_ (.A(_105_),
    .B(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_12.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_115_));
 sky130_fd_sc_hd__xor2_1 _333_ (.A(\CIRCUIT_0.multiply_1.MEMORY_32.s_currentState ),
    .B(_115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_116_));
 sky130_fd_sc_hd__xnor2_1 _334_ (.A(_114_),
    .B(_116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.multiply_1.MEMORY_32.d ));
 sky130_fd_sc_hd__inv_2 _335_ (.A(\CIRCUIT_0.toggle_1.GATES_12.input1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_117_));
 sky130_fd_sc_hd__nor2_1 _336_ (.A(\CIRCUIT_0.toggle_1.GATES_10.input1 ),
    .B(_117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.GATES_10.input1 ));
 sky130_fd_sc_hd__clkbuf_1 _337_ (.A(\CIRCUIT_0.GATES_10.input1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_118_));
 sky130_fd_sc_hd__inv_2 _338_ (.A(_118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_119_));
 sky130_fd_sc_hd__nand4b_1 _339_ (.A_N(\CIRCUIT_0.MEMORY_81.s_currentState ),
    .B(_050_),
    .C(_051_),
    .D(_053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_120_));
 sky130_fd_sc_hd__nor2_2 _340_ (.A(_119_),
    .B(_120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.GATES_59.result ));
 sky130_fd_sc_hd__clkinv_2 _341_ (.A(\CIRCUIT_0.multiply_1.MEMORY_33.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.multiply_1.MEMORY_33.d ));
 sky130_fd_sc_hd__inv_2 _342_ (.A(\CIRCUIT_0.multiply_1.MEMORY_34.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.multiply_1.MEMORY_34.d ));
 sky130_fd_sc_hd__clkbuf_1 _343_ (.A(\CIRCUIT_0.multiply_1.MEMORY_35.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_121_));
 sky130_fd_sc_hd__clkinv_2 _344_ (.A(_121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.multiply_1.GATES_23.input2 ));
 sky130_fd_sc_hd__clkinv_2 _345_ (.A(\CIRCUIT_0.toggle_1.MEMORY_18.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.toggle_1.GATES_10.input2 ));
 sky130_fd_sc_hd__o21bai_1 _346_ (.A1(\CIRCUIT_0.toggle_1.MEMORY_18.s_currentState ),
    .A2(\CIRCUIT_0.toggle_1.GATES_10.input1 ),
    .B1_N(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_122_));
 sky130_fd_sc_hd__a21oi_1 _347_ (.A1(\CIRCUIT_0.toggle_1.MEMORY_18.s_currentState ),
    .A2(_117_),
    .B1(_122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.toggle_1.GATES_12.input1 ));
 sky130_fd_sc_hd__a21oi_1 _348_ (.A1(\CIRCUIT_0.toggle_1.MEMORY_18.s_currentState ),
    .A2(\CIRCUIT_0.toggle_1.GATES_12.input1 ),
    .B1(_122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.toggle_1.GATES_10.input1 ));
 sky130_fd_sc_hd__inv_2 _349_ (.A(\CIRCUIT_0.toggle_1.MEMORY_17.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_123_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _350_ (.A(_123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.output_logic_1.GATES_13.input2 ));
 sky130_fd_sc_hd__clkbuf_1 _351_ (.A(\CIRCUIT_0.inst_dec_1.MEMORY_24.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_124_));
 sky130_fd_sc_hd__clkbuf_1 _352_ (.A(\CIRCUIT_0.inst_dec_1.MEMORY_23.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_125_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _353_ (.A(\CIRCUIT_0.inst_dec_1.MEMORY_22.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_126_));
 sky130_fd_sc_hd__clkbuf_1 _354_ (.A(\CIRCUIT_0.inst_dec_1.MEMORY_21.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_127_));
 sky130_fd_sc_hd__and4b_1 _355_ (.A_N(_124_),
    .B(_125_),
    .C(_126_),
    .D(_127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_128_));
 sky130_fd_sc_hd__clkbuf_1 _356_ (.A(_128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_129_));
 sky130_fd_sc_hd__nor2_1 _357_ (.A(_119_),
    .B(_129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.GATES_65.result ));
 sky130_fd_sc_hd__and2_1 _358_ (.A(\CIRCUIT_0.toggle_1.GATES_10.input1 ),
    .B(_117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_130_));
 sky130_fd_sc_hd__clkbuf_1 _359_ (.A(_130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.dest_reg_sel_1.CLK1 ));
 sky130_fd_sc_hd__or3b_2 _360_ (.A(\CIRCUIT_0.multiply_1.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_0.multiply_1.GATES_24.result ),
    .C_N(clknet_1_1__leaf_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_131_));
 sky130_fd_sc_hd__buf_1 _361_ (.A(_131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_009_));
 sky130_fd_sc_hd__inv_2 _362__1 (.A(clknet_1_1__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net20));
 sky130_fd_sc_hd__inv_2 _362__10 (.A(clknet_1_0__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net29));
 sky130_fd_sc_hd__inv_2 _362__11 (.A(clknet_1_0__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net30));
 sky130_fd_sc_hd__inv_2 _362__12 (.A(clknet_1_0__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net31));
 sky130_fd_sc_hd__inv_2 _362__13 (.A(clknet_1_0__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net32));
 sky130_fd_sc_hd__inv_2 _362__14 (.A(clknet_1_0__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net33));
 sky130_fd_sc_hd__inv_2 _362__15 (.A(clknet_1_1__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net34));
 sky130_fd_sc_hd__inv_2 _362__16 (.A(clknet_1_1__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net35));
 sky130_fd_sc_hd__inv_2 _362__2 (.A(clknet_1_1__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net21));
 sky130_fd_sc_hd__inv_2 _362__3 (.A(clknet_1_1__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net22));
 sky130_fd_sc_hd__inv_2 _362__4 (.A(clknet_1_1__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net23));
 sky130_fd_sc_hd__inv_2 _362__5 (.A(clknet_1_0__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net24));
 sky130_fd_sc_hd__inv_2 _362__6 (.A(clknet_1_1__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net25));
 sky130_fd_sc_hd__inv_2 _362__7 (.A(clknet_1_0__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net26));
 sky130_fd_sc_hd__inv_2 _362__8 (.A(clknet_1_1__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net27));
 sky130_fd_sc_hd__inv_2 _362__9 (.A(clknet_1_0__leaf__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(net28));
 sky130_fd_sc_hd__inv_2 _363_ (.A(\CIRCUIT_0.inst_dec_1.MEMORY_21.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_132_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _364_ (.A(_132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_133_));
 sky130_fd_sc_hd__nor2_1 _365_ (.A(_133_),
    .B(\CIRCUIT_0.MEMORY_76.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_134_));
 sky130_fd_sc_hd__or4_1 _366_ (.A(_127_),
    .B(\CIRCUIT_0.MEMORY_79.s_currentState ),
    .C(\CIRCUIT_0.MEMORY_78.s_currentState ),
    .D(\CIRCUIT_0.MEMORY_77.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_135_));
 sky130_fd_sc_hd__o22a_1 _367_ (.A1(\CIRCUIT_0.inst_dec_1.MEMORY_22.s_currentState ),
    .A2(_134_),
    .B1(_135_),
    .B2(\CIRCUIT_0.MEMORY_75.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_136_));
 sky130_fd_sc_hd__or3b_2 _368_ (.A(_124_),
    .B(_136_),
    .C_N(_125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_137_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _369_ (.A(_137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_138_));
 sky130_fd_sc_hd__mux4_1 _370_ (.A0(\CIRCUIT_0.MEMORY_96.s_currentState ),
    .A1(\CIRCUIT_0.MEMORY_88.s_currentState ),
    .A2(\CIRCUIT_0.MEMORY_77.s_currentState ),
    .A3(_047_),
    .S0(_123_),
    .S1(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_139_));
 sky130_fd_sc_hd__clkbuf_1 _371_ (.A(_139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.O_D0_RR0 ));
 sky130_fd_sc_hd__mux4_1 _372_ (.A0(\CIRCUIT_0.MEMORY_97.s_currentState ),
    .A1(\CIRCUIT_0.MEMORY_89.s_currentState ),
    .A2(_064_),
    .A3(\CIRCUIT_0.MEMORY_81.s_currentState ),
    .S0(_123_),
    .S1(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_140_));
 sky130_fd_sc_hd__clkbuf_1 _373_ (.A(_140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.O_D1_RR1 ));
 sky130_fd_sc_hd__mux4_1 _374_ (.A0(\CIRCUIT_0.MEMORY_98.s_currentState ),
    .A1(\CIRCUIT_0.MEMORY_90.s_currentState ),
    .A2(_059_),
    .A3(\CIRCUIT_0.MEMORY_82.s_currentState ),
    .S0(_123_),
    .S1(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_141_));
 sky130_fd_sc_hd__clkbuf_1 _375_ (.A(_141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.O_D2_RR2 ));
 sky130_fd_sc_hd__mux4_1 _376_ (.A0(\CIRCUIT_0.MEMORY_99.s_currentState ),
    .A1(\CIRCUIT_0.MEMORY_91.s_currentState ),
    .A2(_049_),
    .A3(\CIRCUIT_0.MEMORY_83.s_currentState ),
    .S0(_123_),
    .S1(_137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_142_));
 sky130_fd_sc_hd__clkbuf_1 _377_ (.A(_142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.O_D3_RR3 ));
 sky130_fd_sc_hd__or2_1 _378_ (.A(_124_),
    .B(_125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_143_));
 sky130_fd_sc_hd__clkbuf_1 _379_ (.A(_143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_144_));
 sky130_fd_sc_hd__nand2_1 _380_ (.A(_124_),
    .B(_125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_145_));
 sky130_fd_sc_hd__nand2_1 _381_ (.A(_126_),
    .B(_127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_146_));
 sky130_fd_sc_hd__a21oi_1 _382_ (.A1(_144_),
    .A2(_145_),
    .B1(_146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_147_));
 sky130_fd_sc_hd__mux2_1 _383_ (.A0(\CIRCUIT_0.MEMORY_92.s_currentState ),
    .A1(\CIRCUIT_0.MEMORY_84.s_currentState ),
    .S(_137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_148_));
 sky130_fd_sc_hd__mux2_1 _384_ (.A0(_147_),
    .A1(_148_),
    .S(\CIRCUIT_0.output_logic_1.GATES_13.input2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_149_));
 sky130_fd_sc_hd__clkbuf_1 _385_ (.A(_149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.O_4_MAR ));
 sky130_fd_sc_hd__inv_2 _386_ (.A(_126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_150_));
 sky130_fd_sc_hd__nor2_1 _387_ (.A(\CIRCUIT_0.inst_dec_1.MEMORY_24.s_currentState ),
    .B(\CIRCUIT_0.inst_dec_1.MEMORY_23.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_151_));
 sky130_fd_sc_hd__and4_1 _388_ (.A(_150_),
    .B(_127_),
    .C(_151_),
    .D(_120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_152_));
 sky130_fd_sc_hd__mux2_1 _389_ (.A0(\CIRCUIT_0.MEMORY_93.s_currentState ),
    .A1(\CIRCUIT_0.MEMORY_85.s_currentState ),
    .S(_137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _390_ (.A0(_152_),
    .A1(_153_),
    .S(\CIRCUIT_0.output_logic_1.GATES_13.input2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_154_));
 sky130_fd_sc_hd__clkbuf_1 _391_ (.A(_154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.O_5_WRITE ));
 sky130_fd_sc_hd__o21ba_1 _392_ (.A1(\CIRCUIT_0.toggle_1.MEMORY_17.s_currentState ),
    .A2(\CIRCUIT_0.MEMORY_94.s_currentState ),
    .B1_N(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_155_));
 sky130_fd_sc_hd__a31o_1 _393_ (.A1(\CIRCUIT_0.MEMORY_86.s_currentState ),
    .A2(\CIRCUIT_0.output_logic_1.GATES_13.input2 ),
    .A3(_138_),
    .B1(_155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.O_6_JMP ));
 sky130_fd_sc_hd__mux2_1 _394_ (.A0(\CIRCUIT_0.MEMORY_95.s_currentState ),
    .A1(\CIRCUIT_0.MEMORY_87.s_currentState ),
    .S(_137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_156_));
 sky130_fd_sc_hd__mux2_1 _395_ (.A0(\CIRCUIT_0.MEMORY_74.s_currentState ),
    .A1(_156_),
    .S(\CIRCUIT_0.output_logic_1.GATES_13.input2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_157_));
 sky130_fd_sc_hd__clkbuf_1 _396_ (.A(_157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.O_7_I ));
 sky130_fd_sc_hd__and2b_1 _397_ (.A_N(net16),
    .B(_129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_158_));
 sky130_fd_sc_hd__clkbuf_1 _398_ (.A(_158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.dest_reg_sel_1.GATES_1.result ));
 sky130_fd_sc_hd__nor2_1 _399_ (.A(\CIRCUIT_0.inst_dec_1.MEMORY_22.s_currentState ),
    .B(\CIRCUIT_0.inst_dec_1.MEMORY_21.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_159_));
 sky130_fd_sc_hd__nand2_1 _400_ (.A(_151_),
    .B(_159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_160_));
 sky130_fd_sc_hd__and2_1 _401_ (.A(_049_),
    .B(_160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_161_));
 sky130_fd_sc_hd__xnor2_1 _402_ (.A(_133_),
    .B(_056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_162_));
 sky130_fd_sc_hd__nand2_1 _403_ (.A(_161_),
    .B(_162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_163_));
 sky130_fd_sc_hd__xnor2_1 _404_ (.A(_133_),
    .B(_061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_164_));
 sky130_fd_sc_hd__and2_1 _405_ (.A(_059_),
    .B(_160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_165_));
 sky130_fd_sc_hd__nand2_1 _406_ (.A(_164_),
    .B(_165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_166_));
 sky130_fd_sc_hd__xnor2_1 _407_ (.A(_132_),
    .B(_068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_167_));
 sky130_fd_sc_hd__and2_1 _408_ (.A(_064_),
    .B(_160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_168_));
 sky130_fd_sc_hd__nand2_1 _409_ (.A(_167_),
    .B(_168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_169_));
 sky130_fd_sc_hd__xnor2_1 _410_ (.A(_132_),
    .B(_073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_170_));
 sky130_fd_sc_hd__and2_1 _411_ (.A(\CIRCUIT_0.MEMORY_77.s_currentState ),
    .B(_160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_171_));
 sky130_fd_sc_hd__nand2_1 _412_ (.A(_170_),
    .B(_171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_172_));
 sky130_fd_sc_hd__xor2_1 _413_ (.A(_170_),
    .B(_171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_173_));
 sky130_fd_sc_hd__and3b_1 _414_ (.A_N(\CIRCUIT_0.inst_dec_1.MEMORY_23.s_currentState ),
    .B(\CIRCUIT_0.inst_dec_1.MEMORY_24.s_currentState ),
    .C(\CIRCUIT_0.inst_dec_1.MEMORY_22.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_174_));
 sky130_fd_sc_hd__mux2_1 _415_ (.A0(_127_),
    .A1(\CIRCUIT_0.MEMORY_76.s_currentState ),
    .S(_174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_175_));
 sky130_fd_sc_hd__nand2_1 _416_ (.A(_173_),
    .B(_175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_176_));
 sky130_fd_sc_hd__or2_1 _417_ (.A(_167_),
    .B(_168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_177_));
 sky130_fd_sc_hd__nand2_1 _418_ (.A(_169_),
    .B(_177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_178_));
 sky130_fd_sc_hd__a21o_1 _419_ (.A1(_172_),
    .A2(_176_),
    .B1(_178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_179_));
 sky130_fd_sc_hd__or2_1 _420_ (.A(_164_),
    .B(_165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_180_));
 sky130_fd_sc_hd__nand2_1 _421_ (.A(_166_),
    .B(_180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_181_));
 sky130_fd_sc_hd__a21o_1 _422_ (.A1(_169_),
    .A2(_179_),
    .B1(_181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_182_));
 sky130_fd_sc_hd__xor2_1 _423_ (.A(_161_),
    .B(_162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_183_));
 sky130_fd_sc_hd__inv_2 _424_ (.A(_183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_184_));
 sky130_fd_sc_hd__a21o_1 _425_ (.A1(_166_),
    .A2(_182_),
    .B1(_184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_185_));
 sky130_fd_sc_hd__nand2_1 _426_ (.A(_145_),
    .B(_160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_186_));
 sky130_fd_sc_hd__nand2_1 _427_ (.A(_146_),
    .B(_186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_187_));
 sky130_fd_sc_hd__clkbuf_1 _428_ (.A(_187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_188_));
 sky130_fd_sc_hd__a21boi_1 _429_ (.A1(_163_),
    .A2(_185_),
    .B1_N(_188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.MEMORY_76.d ));
 sky130_fd_sc_hd__clkbuf_1 _430_ (.A(_133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_189_));
 sky130_fd_sc_hd__a21o_1 _431_ (.A1(_159_),
    .A2(_171_),
    .B1(_073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_190_));
 sky130_fd_sc_hd__o211a_1 _432_ (.A1(_189_),
    .A2(\CIRCUIT_0.MEMORY_77.s_currentState ),
    .B1(_190_),
    .C1(_150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_191_));
 sky130_fd_sc_hd__a31o_1 _433_ (.A1(_126_),
    .A2(_189_),
    .A3(_173_),
    .B1(_191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_192_));
 sky130_fd_sc_hd__o21a_1 _434_ (.A1(_173_),
    .A2(_175_),
    .B1(_187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_193_));
 sky130_fd_sc_hd__a32o_1 _435_ (.A1(_146_),
    .A2(_186_),
    .A3(_192_),
    .B1(_193_),
    .B2(_176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.MEMORY_77.d ));
 sky130_fd_sc_hd__nand3_1 _436_ (.A(_178_),
    .B(_172_),
    .C(_176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_194_));
 sky130_fd_sc_hd__nand2_1 _437_ (.A(_126_),
    .B(_189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_195_));
 sky130_fd_sc_hd__nor2_1 _438_ (.A(_178_),
    .B(_195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_196_));
 sky130_fd_sc_hd__and3_1 _439_ (.A(_064_),
    .B(_144_),
    .C(_159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_197_));
 sky130_fd_sc_hd__o221a_1 _440_ (.A1(_189_),
    .A2(_064_),
    .B1(_068_),
    .B2(_197_),
    .C1(_150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_198_));
 sky130_fd_sc_hd__o21ba_1 _441_ (.A1(_196_),
    .A2(_198_),
    .B1_N(_187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_199_));
 sky130_fd_sc_hd__a31o_1 _442_ (.A1(_179_),
    .A2(_188_),
    .A3(_194_),
    .B1(_199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.MEMORY_78.d ));
 sky130_fd_sc_hd__nand3_1 _443_ (.A(_181_),
    .B(_169_),
    .C(_179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_200_));
 sky130_fd_sc_hd__and3_1 _444_ (.A(_059_),
    .B(_144_),
    .C(_159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_201_));
 sky130_fd_sc_hd__o221a_1 _445_ (.A1(_189_),
    .A2(_059_),
    .B1(_061_),
    .B2(_201_),
    .C1(_150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_202_));
 sky130_fd_sc_hd__o21ba_1 _446_ (.A1(_181_),
    .A2(_195_),
    .B1_N(_202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_203_));
 sky130_fd_sc_hd__nor2_1 _447_ (.A(_187_),
    .B(_203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_204_));
 sky130_fd_sc_hd__a31o_1 _448_ (.A1(_182_),
    .A2(_188_),
    .A3(_200_),
    .B1(_204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.MEMORY_79.d ));
 sky130_fd_sc_hd__nand3_1 _449_ (.A(_184_),
    .B(_166_),
    .C(_182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_205_));
 sky130_fd_sc_hd__and3_1 _450_ (.A(_049_),
    .B(_143_),
    .C(_159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_206_));
 sky130_fd_sc_hd__o221a_1 _451_ (.A1(_049_),
    .A2(_133_),
    .B1(_056_),
    .B2(_206_),
    .C1(_150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_207_));
 sky130_fd_sc_hd__o21ba_1 _452_ (.A1(_184_),
    .A2(_195_),
    .B1_N(_207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_208_));
 sky130_fd_sc_hd__nor2_1 _453_ (.A(_187_),
    .B(_208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_209_));
 sky130_fd_sc_hd__a31o_1 _454_ (.A1(_185_),
    .A2(_188_),
    .A3(_205_),
    .B1(_209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.MEMORY_75.d ));
 sky130_fd_sc_hd__or2_1 _455_ (.A(_118_),
    .B(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_210_));
 sky130_fd_sc_hd__clkbuf_1 _456_ (.A(_210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.toggle_1.GATES_8.result ));
 sky130_fd_sc_hd__nor2_1 _457_ (.A(_144_),
    .B(_195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.MEMORY_74.d ));
 sky130_fd_sc_hd__o21a_1 _458_ (.A1(_119_),
    .A2(_129_),
    .B1(\CIRCUIT_0.MEMORY_100.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.GATES_72.result ));
 sky130_fd_sc_hd__and3_1 _459_ (.A(\CIRCUIT_0.dest_reg_sel_1.MEMORY_2.s_currentState ),
    .B(_118_),
    .C(_129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_211_));
 sky130_fd_sc_hd__clkbuf_1 _460_ (.A(_211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.GATES_43.result ));
 sky130_fd_sc_hd__nor3_1 _461_ (.A(net16),
    .B(_146_),
    .C(_145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.GATES_42.result ));
 sky130_fd_sc_hd__and3_1 _462_ (.A(\CIRCUIT_0.dest_reg_sel_1.MEMORY_4.s_currentState ),
    .B(_118_),
    .C(_129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_212_));
 sky130_fd_sc_hd__clkbuf_1 _463_ (.A(_212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.GATES_41.result ));
 sky130_fd_sc_hd__and3_1 _464_ (.A(\CIRCUIT_0.dest_reg_sel_1.MEMORY_3.s_currentState ),
    .B(_118_),
    .C(_128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_213_));
 sky130_fd_sc_hd__clkbuf_1 _465_ (.A(_213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.GATES_40.result ));
 sky130_fd_sc_hd__nor3_1 _466_ (.A(net16),
    .B(_144_),
    .C(_146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.GATES_39.result ));
 sky130_fd_sc_hd__and3b_1 _467_ (.A_N(_125_),
    .B(\CIRCUIT_0.GATES_10.input1 ),
    .C(_124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_214_));
 sky130_fd_sc_hd__clkbuf_1 _468_ (.A(_214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\CIRCUIT_0.GATES_11.result ));
 sky130_fd_sc_hd__o21bai_1 _469_ (.A1(_119_),
    .A2(_188_),
    .B1_N(\CIRCUIT_0.GATES_11.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.GATES_10.result ));
 sky130_fd_sc_hd__a21oi_1 _470_ (.A1(_105_),
    .A2(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_13.s_currentState ),
    .B1(\CIRCUIT_0.multiply_1.MEMORY_25.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_215_));
 sky130_fd_sc_hd__nor2_1 _471_ (.A(_086_),
    .B(_215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.multiply_1.MEMORY_25.d ));
 sky130_fd_sc_hd__a21oi_1 _472_ (.A1(_085_),
    .A2(_087_),
    .B1(_086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_216_));
 sky130_fd_sc_hd__nor2_1 _473_ (.A(_088_),
    .B(_216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\CIRCUIT_0.multiply_1.MEMORY_26.d ));
 sky130_fd_sc_hd__clkbuf_2 _474_ (.A(\CIRCUIT_0.GATES_59.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_217_));
 sky130_fd_sc_hd__inv_2 _475_ (.A(_217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _476_ (.A(_217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _477_ (.A(_217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _478_ (.A(_217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _479_ (.A(_217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _480_ (.A(\CIRCUIT_0.GATES_59.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _481_ (.A(\CIRCUIT_0.GATES_59.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _482_ (.A(\CIRCUIT_0.multiply_1.MEMORY_33.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_011_));
 sky130_fd_sc_hd__clkinv_2 _483_ (.A(\CIRCUIT_0.multiply_1.MEMORY_34.s_currentState ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_013_));
 sky130_fd_sc_hd__nand2_1 _484_ (.A(_083_),
    .B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_015_));
 sky130_fd_sc_hd__nand2_1 _485_ (.A(_083_),
    .B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_017_));
 sky130_fd_sc_hd__nand2_1 _486_ (.A(_083_),
    .B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_019_));
 sky130_fd_sc_hd__nand2_1 _487_ (.A(_083_),
    .B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_021_));
 sky130_fd_sc_hd__buf_1 _488_ (.A(clknet_1_1__leaf_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_218_));
 sky130_fd_sc_hd__or3b_2 _489_ (.A(_121_),
    .B(_077_),
    .C_N(clknet_1_0__leaf__218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_219_));
 sky130_fd_sc_hd__buf_1 _490_ (.A(_219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_023_));
 sky130_fd_sc_hd__or3b_2 _491_ (.A(_121_),
    .B(_077_),
    .C_N(clknet_1_1__leaf__218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_220_));
 sky130_fd_sc_hd__buf_1 _492_ (.A(_220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_025_));
 sky130_fd_sc_hd__or3b_2 _493_ (.A(_121_),
    .B(_077_),
    .C_N(clknet_1_0__leaf__218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_221_));
 sky130_fd_sc_hd__buf_1 _494_ (.A(_221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_027_));
 sky130_fd_sc_hd__or3b_2 _495_ (.A(_121_),
    .B(\CIRCUIT_0.multiply_1.GATES_24.result ),
    .C_N(clknet_1_1__leaf__218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_222_));
 sky130_fd_sc_hd__buf_1 _496_ (.A(_222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_029_));
 sky130_fd_sc_hd__nor2_1 _497_ (.A(_047_),
    .B(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_223_));
 sky130_fd_sc_hd__nand2_1 _498_ (.A(_223_),
    .B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_031_));
 sky130_fd_sc_hd__nand2_1 _499_ (.A(_223_),
    .B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_033_));
 sky130_fd_sc_hd__nand2_1 _500_ (.A(_223_),
    .B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_035_));
 sky130_fd_sc_hd__nand2_1 _501_ (.A(_223_),
    .B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_037_));
 sky130_fd_sc_hd__clkbuf_2 _502_ (.A(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_224_));
 sky130_fd_sc_hd__clkbuf_2 _503_ (.A(_224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_225_));
 sky130_fd_sc_hd__buf_1 _504_ (.A(clknet_1_1__leaf__218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_226_));
 sky130_fd_sc_hd__buf_1 _505_ (.A(clknet_1_1__leaf__226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_227_));
 sky130_fd_sc_hd__nand2_2 _506_ (.A(_225_),
    .B(clknet_1_1__leaf__227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_038_));
 sky130_fd_sc_hd__nand2_2 _507_ (.A(_225_),
    .B(clknet_1_0__leaf__227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_039_));
 sky130_fd_sc_hd__nand2_2 _508_ (.A(_225_),
    .B(clknet_1_1__leaf__227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_040_));
 sky130_fd_sc_hd__nand2_2 _509_ (.A(_225_),
    .B(clknet_1_1__leaf__227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_041_));
 sky130_fd_sc_hd__nand2_2 _510_ (.A(_225_),
    .B(clknet_1_0__leaf__227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_042_));
 sky130_fd_sc_hd__nand2_2 _511_ (.A(_224_),
    .B(clknet_1_0__leaf__226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_043_));
 sky130_fd_sc_hd__nand2_2 _512_ (.A(_224_),
    .B(clknet_1_0__leaf__226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_044_));
 sky130_fd_sc_hd__nand2_2 _513_ (.A(_224_),
    .B(clknet_1_0__leaf__226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_045_));
 sky130_fd_sc_hd__nand2_2 _514_ (.A(_224_),
    .B(clknet_1_0__leaf__226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_046_));
 sky130_fd_sc_hd__dfrtp_1 _515_ (.CLK(net35),
    .D(\CIRCUIT_0.multiply_1.MEMORY_25.d ),
    .RESET_B(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_25.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _516_ (.CLK(net34),
    .D(\CIRCUIT_0.multiply_1.MEMORY_26.d ),
    .RESET_B(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_26.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _517_ (.CLK(net33),
    .D(\CIRCUIT_0.multiply_1.MEMORY_27.d ),
    .RESET_B(_002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_27.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _518_ (.CLK(net32),
    .D(\CIRCUIT_0.multiply_1.MEMORY_28.d ),
    .RESET_B(_003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_28.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _519_ (.CLK(net31),
    .D(\CIRCUIT_0.multiply_1.MEMORY_29.d ),
    .RESET_B(_004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_29.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _520_ (.CLK(net30),
    .D(\CIRCUIT_0.multiply_1.MEMORY_30.d ),
    .RESET_B(_005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_30.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _521_ (.CLK(net29),
    .D(\CIRCUIT_0.multiply_1.MEMORY_31.d ),
    .RESET_B(_006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_31.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _522_ (.CLK(net28),
    .D(\CIRCUIT_0.multiply_1.MEMORY_32.d ),
    .RESET_B(_007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_32.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _523_ (.CLK(clknet_1_0__leaf__009_),
    .D(\CIRCUIT_0.multiply_1.MEMORY_33.d ),
    .RESET_B(_008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_33.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _524_ (.CLK(_011_),
    .D(\CIRCUIT_0.multiply_1.MEMORY_34.d ),
    .RESET_B(_010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_34.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _525_ (.CLK(_013_),
    .D(\CIRCUIT_0.multiply_1.GATES_23.input2 ),
    .RESET_B(_012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.MEMORY_35.s_currentState ));
 sky130_fd_sc_hd__dfbbn_1 _526_ (.CLK_N(net27),
    .D(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_15.s_currentState ),
    .RESET_B(_014_),
    .SET_B(_015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_16.s_currentState ),
    .Q_N(_235_));
 sky130_fd_sc_hd__dfbbn_1 _527_ (.CLK_N(net26),
    .D(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_14.s_currentState ),
    .RESET_B(_016_),
    .SET_B(_017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_15.s_currentState ),
    .Q_N(_234_));
 sky130_fd_sc_hd__dfbbn_1 _528_ (.CLK_N(net25),
    .D(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_13.s_currentState ),
    .RESET_B(_018_),
    .SET_B(_019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_14.s_currentState ),
    .Q_N(_233_));
 sky130_fd_sc_hd__dfbbn_1 _529_ (.CLK_N(net24),
    .D(net18),
    .RESET_B(_020_),
    .SET_B(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_13.s_currentState ),
    .Q_N(_232_));
 sky130_fd_sc_hd__conb_1 _529__18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net18));
 sky130_fd_sc_hd__dfrtp_1 _530_ (.CLK(_023_),
    .D(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_11.s_currentState ),
    .RESET_B(_022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_12.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _531_ (.CLK(_025_),
    .D(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_10.s_currentState ),
    .RESET_B(_024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_11.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _532_ (.CLK(_027_),
    .D(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_9.s_currentState ),
    .RESET_B(_026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_10.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _533_ (.CLK(_029_),
    .D(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_16.s_currentState ),
    .RESET_B(_028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_8_1.MEMORY_9.s_currentState ));
 sky130_fd_sc_hd__dfbbn_1 _534_ (.CLK_N(net23),
    .D(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_11.s_currentState ),
    .RESET_B(_030_),
    .SET_B(_031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_12.s_currentState ),
    .Q_N(_231_));
 sky130_fd_sc_hd__dfbbn_1 _535_ (.CLK_N(net22),
    .D(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_10.s_currentState ),
    .RESET_B(_032_),
    .SET_B(_033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_11.s_currentState ),
    .Q_N(_230_));
 sky130_fd_sc_hd__dfbbn_1 _536_ (.CLK_N(net21),
    .D(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_9.s_currentState ),
    .RESET_B(_034_),
    .SET_B(_035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_10.s_currentState ),
    .Q_N(_229_));
 sky130_fd_sc_hd__dfbbn_1 _537_ (.CLK_N(net20),
    .D(net19),
    .RESET_B(_036_),
    .SET_B(_037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.multiply_1.shift_reg_1.MEMORY_9.s_currentState ),
    .Q_N(_228_));
 sky130_fd_sc_hd__conb_1 _537__19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net19));
 sky130_fd_sc_hd__dfstp_1 _538_ (.CLK(\CIRCUIT_0.dest_reg_sel_1.GATES_1.result ),
    .D(\CIRCUIT_0.dest_reg_sel_1.MEMORY_4.s_currentState ),
    .SET_B(_038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.dest_reg_sel_1.MEMORY_2.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _539_ (.CLK(\CIRCUIT_0.dest_reg_sel_1.GATES_1.result ),
    .D(\CIRCUIT_0.dest_reg_sel_1.MEMORY_2.s_currentState ),
    .RESET_B(_039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.dest_reg_sel_1.MEMORY_3.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _540_ (.CLK(\CIRCUIT_0.dest_reg_sel_1.GATES_1.result ),
    .D(\CIRCUIT_0.dest_reg_sel_1.MEMORY_3.s_currentState ),
    .RESET_B(_040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.dest_reg_sel_1.MEMORY_4.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _541_ (.CLK(\CIRCUIT_0.toggle_1.GATES_8.result ),
    .D(\CIRCUIT_0.output_logic_1.GATES_13.input2 ),
    .SET_B(_041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.toggle_1.MEMORY_17.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _542_ (.CLK(clknet_1_0__leaf_io_in[0]),
    .D(\CIRCUIT_0.toggle_1.GATES_10.input2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.toggle_1.MEMORY_18.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _543_ (.CLK(\CIRCUIT_0.dest_reg_sel_1.CLK1 ),
    .D(net2),
    .RESET_B(_042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.inst_dec_1.MEMORY_21.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _544_ (.CLK(net17),
    .D(net3),
    .RESET_B(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.inst_dec_1.MEMORY_22.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _545_ (.CLK(net17),
    .D(net4),
    .RESET_B(_044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.inst_dec_1.MEMORY_23.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _546_ (.CLK(net17),
    .D(net5),
    .RESET_B(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.inst_dec_1.MEMORY_24.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _547_ (.CLK(clknet_1_0__leaf_io_in[0]),
    .D(\CIRCUIT_0.GATES_65.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_100.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _548_ (.CLK(\CIRCUIT_0.GATES_43.result ),
    .D(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_99.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _549_ (.CLK(\CIRCUIT_0.GATES_43.result ),
    .D(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_98.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _550_ (.CLK(\CIRCUIT_0.GATES_43.result ),
    .D(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_97.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _551_ (.CLK(\CIRCUIT_0.GATES_43.result ),
    .D(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_96.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _552_ (.CLK(\CIRCUIT_0.GATES_41.result ),
    .D(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_95.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _553_ (.CLK(\CIRCUIT_0.GATES_41.result ),
    .D(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_94.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _554_ (.CLK(\CIRCUIT_0.GATES_41.result ),
    .D(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_93.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _555_ (.CLK(\CIRCUIT_0.GATES_41.result ),
    .D(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_92.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _556_ (.CLK(\CIRCUIT_0.GATES_40.result ),
    .D(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_91.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _557_ (.CLK(\CIRCUIT_0.GATES_40.result ),
    .D(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_90.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _558_ (.CLK(\CIRCUIT_0.GATES_40.result ),
    .D(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_89.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _559_ (.CLK(\CIRCUIT_0.GATES_40.result ),
    .D(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_88.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _560_ (.CLK(\CIRCUIT_0.GATES_42.result ),
    .D(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_87.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _561_ (.CLK(\CIRCUIT_0.GATES_42.result ),
    .D(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_86.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _562_ (.CLK(\CIRCUIT_0.GATES_42.result ),
    .D(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_85.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _563_ (.CLK(\CIRCUIT_0.GATES_42.result ),
    .D(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_84.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _564_ (.CLK(\CIRCUIT_0.GATES_39.result ),
    .D(\CIRCUIT_0.GATES_36.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_83.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _565_ (.CLK(\CIRCUIT_0.GATES_39.result ),
    .D(\CIRCUIT_0.GATES_31.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_82.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _566_ (.CLK(\CIRCUIT_0.GATES_39.result ),
    .D(\CIRCUIT_0.GATES_29.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_81.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _567_ (.CLK(\CIRCUIT_0.GATES_39.result ),
    .D(\CIRCUIT_0.GATES_28.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_80.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _568_ (.CLK(\CIRCUIT_0.GATES_10.result ),
    .D(\CIRCUIT_0.MEMORY_79.d ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_79.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _569_ (.CLK(\CIRCUIT_0.GATES_10.result ),
    .D(\CIRCUIT_0.MEMORY_78.d ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_78.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _570_ (.CLK(\CIRCUIT_0.GATES_10.result ),
    .D(\CIRCUIT_0.MEMORY_77.d ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_77.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _571_ (.CLK(\CIRCUIT_0.GATES_11.result ),
    .D(\CIRCUIT_0.MEMORY_76.d ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_76.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _572_ (.CLK(\CIRCUIT_0.GATES_10.result ),
    .D(\CIRCUIT_0.MEMORY_75.d ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_75.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _573_ (.CLK(\CIRCUIT_0.GATES_72.result ),
    .D(\CIRCUIT_0.MEMORY_74.d ),
    .RESET_B(_046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\CIRCUIT_0.MEMORY_74.s_currentState ));
 sky130_fd_sc_hd__buf_2 _576_ (.A(\CIRCUIT_0.O_D0_RR0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 _577_ (.A(\CIRCUIT_0.O_D1_RR1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_2 _578_ (.A(\CIRCUIT_0.O_D2_RR2 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_2 _579_ (.A(\CIRCUIT_0.O_D3_RR3 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_2 _580_ (.A(\CIRCUIT_0.O_4_MAR ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 _581_ (.A(\CIRCUIT_0.O_5_WRITE ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 _582_ (.A(\CIRCUIT_0.O_6_JMP ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 _583_ (.A(\CIRCUIT_0.O_7_I ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__009_ (.A(_009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0__009_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__218_ (.A(_218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0__218_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__226_ (.A(_226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0__226_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__227_ (.A(_227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0__227_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_io_in[0]  (.A(io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__009_ (.A(clknet_0__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_0__leaf__009_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__218_ (.A(clknet_0__218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_0__leaf__218_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__226_ (.A(clknet_0__226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_0__leaf__226_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__227_ (.A(clknet_0__227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_0__leaf__227_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_0__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__009_ (.A(clknet_0__009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_1__leaf__009_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__218_ (.A(clknet_0__218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_1__leaf__218_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__226_ (.A(clknet_0__226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_1__leaf__226_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__227_ (.A(clknet_0__227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_1__leaf__227_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_1__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(io_in[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(io_in[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 repeater10 (.A(\CIRCUIT_0.GATES_29.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 repeater11 (.A(\CIRCUIT_0.GATES_29.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 repeater12 (.A(\CIRCUIT_0.GATES_31.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 repeater13 (.A(\CIRCUIT_0.GATES_31.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 repeater14 (.A(\CIRCUIT_0.GATES_36.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 repeater15 (.A(\CIRCUIT_0.GATES_36.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 repeater16 (.A(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 repeater17 (.A(\CIRCUIT_0.dest_reg_sel_1.CLK1 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 repeater8 (.A(\CIRCUIT_0.GATES_28.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 repeater9 (.A(\CIRCUIT_0.GATES_28.result ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net9));
endmodule
