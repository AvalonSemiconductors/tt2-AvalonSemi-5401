magic
tech sky130A
magscale 1 2
timestamp 1667177659
<< obsli1 >>
rect 1104 1071 16836 22865
<< obsm1 >>
rect 1104 1040 16836 22896
<< obsm2 >>
rect 1306 711 15076 23225
<< metal3 >>
rect 0 23128 400 23248
rect 0 21632 400 21752
rect 0 20136 400 20256
rect 0 18640 400 18760
rect 0 17144 400 17264
rect 0 15648 400 15768
rect 0 14152 400 14272
rect 0 12656 400 12776
rect 0 11160 400 11280
rect 0 9664 400 9784
rect 0 8168 400 8288
rect 0 6672 400 6792
rect 0 5176 400 5296
rect 0 3680 400 3800
rect 0 2184 400 2304
rect 0 688 400 808
<< obsm3 >>
rect 480 23048 15080 23221
rect 400 21832 15080 23048
rect 480 21552 15080 21832
rect 400 20336 15080 21552
rect 480 20056 15080 20336
rect 400 18840 15080 20056
rect 480 18560 15080 18840
rect 400 17344 15080 18560
rect 480 17064 15080 17344
rect 400 15848 15080 17064
rect 480 15568 15080 15848
rect 400 14352 15080 15568
rect 480 14072 15080 14352
rect 400 12856 15080 14072
rect 480 12576 15080 12856
rect 400 11360 15080 12576
rect 480 11080 15080 11360
rect 400 9864 15080 11080
rect 480 9584 15080 9864
rect 400 8368 15080 9584
rect 480 8088 15080 8368
rect 400 6872 15080 8088
rect 480 6592 15080 6872
rect 400 5376 15080 6592
rect 480 5096 15080 5376
rect 400 3880 15080 5096
rect 480 3600 15080 3880
rect 400 2384 15080 3600
rect 480 2104 15080 2384
rect 400 888 15080 2104
rect 480 715 15080 888
<< metal4 >>
rect 2918 1040 3238 22896
rect 4892 1040 5212 22896
rect 6866 1040 7186 22896
rect 8840 1040 9160 22896
rect 10814 1040 11134 22896
rect 12788 1040 13108 22896
rect 14762 1040 15082 22896
<< obsm4 >>
rect 2635 3027 2838 15469
rect 3318 3027 4812 15469
rect 5292 3027 6786 15469
rect 7266 3027 8760 15469
rect 9240 3027 10734 15469
rect 11214 3027 11349 15469
<< labels >>
rlabel metal3 s 0 688 400 808 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 2184 400 2304 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 0 3680 400 3800 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 0 5176 400 5296 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 0 6672 400 6792 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 0 8168 400 8288 6 io_in[5]
port 6 nsew signal input
rlabel metal3 s 0 9664 400 9784 6 io_in[6]
port 7 nsew signal input
rlabel metal3 s 0 11160 400 11280 6 io_in[7]
port 8 nsew signal input
rlabel metal3 s 0 12656 400 12776 6 io_out[0]
port 9 nsew signal output
rlabel metal3 s 0 14152 400 14272 6 io_out[1]
port 10 nsew signal output
rlabel metal3 s 0 15648 400 15768 6 io_out[2]
port 11 nsew signal output
rlabel metal3 s 0 17144 400 17264 6 io_out[3]
port 12 nsew signal output
rlabel metal3 s 0 18640 400 18760 6 io_out[4]
port 13 nsew signal output
rlabel metal3 s 0 20136 400 20256 6 io_out[5]
port 14 nsew signal output
rlabel metal3 s 0 21632 400 21752 6 io_out[6]
port 15 nsew signal output
rlabel metal3 s 0 23128 400 23248 6 io_out[7]
port 16 nsew signal output
rlabel metal4 s 2918 1040 3238 22896 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 6866 1040 7186 22896 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 10814 1040 11134 22896 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 14762 1040 15082 22896 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 4892 1040 5212 22896 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 8840 1040 9160 22896 6 vssd1
port 18 nsew ground bidirectional
rlabel metal4 s 12788 1040 13108 22896 6 vssd1
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 18000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1079892
string GDS_FILE /work/runs/wokwi/results/signoff/tholin_avalonsemi_5401.magic.gds
string GDS_START 290208
<< end >>

