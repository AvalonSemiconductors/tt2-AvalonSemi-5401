magic
tech sky130A
magscale 1 2
timestamp 1668080783
<< checkpaint >>
rect -3932 -3930 21675 27180
<< viali >>
rect 1409 22593 1443 22627
rect 1593 22593 1627 22627
rect 1501 22457 1535 22491
rect 1961 22389 1995 22423
rect 1593 22185 1627 22219
rect 2789 22117 2823 22151
rect 1409 21981 1443 22015
rect 2329 21981 2363 22015
rect 2973 21981 3007 22015
rect 2145 21845 2179 21879
rect 1501 21505 1535 21539
rect 2237 21505 2271 21539
rect 3157 21505 3191 21539
rect 3801 21505 3835 21539
rect 2973 21369 3007 21403
rect 1685 21301 1719 21335
rect 2421 21301 2455 21335
rect 3617 21301 3651 21335
rect 2421 21097 2455 21131
rect 1501 20893 1535 20927
rect 2237 20893 2271 20927
rect 2973 20893 3007 20927
rect 3985 20893 4019 20927
rect 4629 20893 4663 20927
rect 1685 20757 1719 20791
rect 3157 20757 3191 20791
rect 3801 20757 3835 20791
rect 4445 20757 4479 20791
rect 3709 20553 3743 20587
rect 4077 20553 4111 20587
rect 4905 20553 4939 20587
rect 1593 20417 1627 20451
rect 2053 20417 2087 20451
rect 2789 20417 2823 20451
rect 3525 20417 3559 20451
rect 4261 20417 4295 20451
rect 5089 20417 5123 20451
rect 5733 20417 5767 20451
rect 3065 20349 3099 20383
rect 4629 20349 4663 20383
rect 2789 20281 2823 20315
rect 2881 20281 2915 20315
rect 1409 20213 1443 20247
rect 2237 20213 2271 20247
rect 5549 20213 5583 20247
rect 2421 20009 2455 20043
rect 3065 19941 3099 19975
rect 3801 19941 3835 19975
rect 5365 19941 5399 19975
rect 1777 19873 1811 19907
rect 2145 19805 2179 19839
rect 2237 19805 2271 19839
rect 2973 19805 3007 19839
rect 3249 19805 3283 19839
rect 3985 19805 4019 19839
rect 4077 19805 4111 19839
rect 4537 19805 4571 19839
rect 5181 19805 5215 19839
rect 5825 19805 5859 19839
rect 6021 19805 6055 19839
rect 6653 19805 6687 19839
rect 3801 19737 3835 19771
rect 5917 19737 5951 19771
rect 2973 19669 3007 19703
rect 4629 19669 4663 19703
rect 6469 19669 6503 19703
rect 1409 19465 1443 19499
rect 3725 19465 3759 19499
rect 7113 19465 7147 19499
rect 3525 19397 3559 19431
rect 4905 19397 4939 19431
rect 6469 19397 6503 19431
rect 5135 19363 5169 19397
rect 1593 19329 1627 19363
rect 1685 19329 1719 19363
rect 1961 19329 1995 19363
rect 2789 19329 2823 19363
rect 2973 19329 3007 19363
rect 6377 19329 6411 19363
rect 6561 19329 6595 19363
rect 7021 19329 7055 19363
rect 2053 19261 2087 19295
rect 3065 19261 3099 19295
rect 3893 19193 3927 19227
rect 3709 19125 3743 19159
rect 5089 19125 5123 19159
rect 5273 19125 5307 19159
rect 2513 18921 2547 18955
rect 7205 18921 7239 18955
rect 4261 18853 4295 18887
rect 7757 18853 7791 18887
rect 3065 18785 3099 18819
rect 1685 18717 1719 18751
rect 1869 18717 1903 18751
rect 5457 18717 5491 18751
rect 5733 18717 5767 18751
rect 6193 18717 6227 18751
rect 6469 18717 6503 18751
rect 6561 18717 6595 18751
rect 7113 18717 7147 18751
rect 7941 18717 7975 18751
rect 1961 18649 1995 18683
rect 3985 18649 4019 18683
rect 5273 18649 5307 18683
rect 2881 18581 2915 18615
rect 2973 18581 3007 18615
rect 4445 18581 4479 18615
rect 5641 18581 5675 18615
rect 6561 18377 6595 18411
rect 7481 18377 7515 18411
rect 8677 18377 8711 18411
rect 9505 18377 9539 18411
rect 6377 18309 6411 18343
rect 8125 18309 8159 18343
rect 2125 18241 2159 18275
rect 4057 18241 4091 18275
rect 5641 18241 5675 18275
rect 7389 18241 7423 18275
rect 8033 18241 8067 18275
rect 8217 18241 8251 18275
rect 8861 18241 8895 18275
rect 9321 18241 9355 18275
rect 9505 18241 9539 18275
rect 1869 18173 1903 18207
rect 3801 18173 3835 18207
rect 5825 18105 5859 18139
rect 6745 18105 6779 18139
rect 3249 18037 3283 18071
rect 5181 18037 5215 18071
rect 6561 18037 6595 18071
rect 5641 17833 5675 17867
rect 6377 17833 6411 17867
rect 8953 17833 8987 17867
rect 3249 17765 3283 17799
rect 8217 17765 8251 17799
rect 1869 17629 1903 17663
rect 4261 17629 4295 17663
rect 6653 17629 6687 17663
rect 7297 17629 7331 17663
rect 7573 17629 7607 17663
rect 8217 17629 8251 17663
rect 8401 17629 8435 17663
rect 9137 17629 9171 17663
rect 9597 17629 9631 17663
rect 9789 17629 9823 17663
rect 2114 17561 2148 17595
rect 4506 17561 4540 17595
rect 6193 17561 6227 17595
rect 7113 17561 7147 17595
rect 7481 17561 7515 17595
rect 6377 17493 6411 17527
rect 9781 17493 9815 17527
rect 3341 17289 3375 17323
rect 4046 17221 4080 17255
rect 7757 17221 7791 17255
rect 1961 17153 1995 17187
rect 2228 17153 2262 17187
rect 3801 17153 3835 17187
rect 5825 17153 5859 17187
rect 6561 17153 6595 17187
rect 6653 17153 6687 17187
rect 6837 17153 6871 17187
rect 7573 17153 7607 17187
rect 7849 17153 7883 17187
rect 8401 17153 8435 17187
rect 9045 17153 9079 17187
rect 9689 17153 9723 17187
rect 9873 17153 9907 17187
rect 10517 17153 10551 17187
rect 7389 17085 7423 17119
rect 5641 17017 5675 17051
rect 6745 17017 6779 17051
rect 10149 17017 10183 17051
rect 10701 17017 10735 17051
rect 5181 16949 5215 16983
rect 6377 16949 6411 16983
rect 8493 16949 8527 16983
rect 9137 16949 9171 16983
rect 9781 16949 9815 16983
rect 6561 16745 6595 16779
rect 10609 16745 10643 16779
rect 11529 16677 11563 16711
rect 1869 16541 1903 16575
rect 4537 16541 4571 16575
rect 7941 16541 7975 16575
rect 8125 16541 8159 16575
rect 8401 16541 8435 16575
rect 11713 16541 11747 16575
rect 2114 16473 2148 16507
rect 4261 16473 4295 16507
rect 5273 16473 5307 16507
rect 9321 16473 9355 16507
rect 3249 16405 3283 16439
rect 4445 16405 4479 16439
rect 4629 16405 4663 16439
rect 4813 16405 4847 16439
rect 8309 16405 8343 16439
rect 1409 16201 1443 16235
rect 15301 16201 15335 16235
rect 2872 16133 2906 16167
rect 4712 16133 4746 16167
rect 6929 16133 6963 16167
rect 8213 16133 8247 16167
rect 10793 16133 10827 16167
rect 1685 16065 1719 16099
rect 1777 16065 1811 16099
rect 6377 16065 6411 16099
rect 6653 16065 6687 16099
rect 7205 16065 7239 16099
rect 7941 16065 7975 16099
rect 8125 16065 8159 16099
rect 8309 16065 8343 16099
rect 9689 16065 9723 16099
rect 9873 16065 9907 16099
rect 9965 16065 9999 16099
rect 10609 16065 10643 16099
rect 10885 16065 10919 16099
rect 11713 16065 11747 16099
rect 12357 16065 12391 16099
rect 15485 16065 15519 16099
rect 1593 15997 1627 16031
rect 1869 15997 1903 16031
rect 2605 15997 2639 16031
rect 4445 15997 4479 16031
rect 3985 15861 4019 15895
rect 5825 15861 5859 15895
rect 8493 15861 8527 15895
rect 9505 15861 9539 15895
rect 10425 15861 10459 15895
rect 11529 15861 11563 15895
rect 12173 15861 12207 15895
rect 3985 15657 4019 15691
rect 4813 15657 4847 15691
rect 6561 15657 6595 15691
rect 13093 15657 13127 15691
rect 14565 15657 14599 15691
rect 10931 15589 10965 15623
rect 12357 15589 12391 15623
rect 8125 15521 8159 15555
rect 11069 15521 11103 15555
rect 11161 15521 11195 15555
rect 1409 15453 1443 15487
rect 3985 15453 4019 15487
rect 4169 15453 4203 15487
rect 4629 15453 4663 15487
rect 5273 15453 5307 15487
rect 7849 15453 7883 15487
rect 9156 15453 9190 15487
rect 9413 15453 9447 15487
rect 10057 15453 10091 15487
rect 10241 15453 10275 15487
rect 10333 15453 10367 15487
rect 10793 15453 10827 15487
rect 11253 15453 11287 15487
rect 11713 15453 11747 15487
rect 11897 15453 11931 15487
rect 12541 15453 12575 15487
rect 13001 15453 13035 15487
rect 13185 15453 13219 15487
rect 14381 15453 14415 15487
rect 15577 15453 15611 15487
rect 1654 15385 1688 15419
rect 2789 15317 2823 15351
rect 7481 15317 7515 15351
rect 7941 15317 7975 15351
rect 8953 15317 8987 15351
rect 9321 15317 9355 15351
rect 9873 15317 9907 15351
rect 11805 15317 11839 15351
rect 15761 15317 15795 15351
rect 1409 15113 1443 15147
rect 11713 15113 11747 15147
rect 13829 15113 13863 15147
rect 15669 15113 15703 15147
rect 4690 15045 4724 15079
rect 6929 15045 6963 15079
rect 8033 15045 8067 15079
rect 10425 15045 10459 15079
rect 11529 15045 11563 15079
rect 1602 14977 1636 15011
rect 1869 14977 1903 15011
rect 2053 14977 2087 15011
rect 2872 14977 2906 15011
rect 6469 14977 6503 15011
rect 6653 14977 6687 15011
rect 7205 14977 7239 15011
rect 10241 14977 10275 15011
rect 10517 14977 10551 15011
rect 10609 14977 10643 15011
rect 11989 14977 12023 15011
rect 12441 14977 12475 15011
rect 13093 14977 13127 15011
rect 13737 14977 13771 15011
rect 14933 14977 14967 15011
rect 15577 14977 15611 15011
rect 2605 14909 2639 14943
rect 4445 14909 4479 14943
rect 12633 14841 12667 14875
rect 15117 14841 15151 14875
rect 3985 14773 4019 14807
rect 5825 14773 5859 14807
rect 9321 14773 9355 14807
rect 10793 14773 10827 14807
rect 11713 14773 11747 14807
rect 13277 14773 13311 14807
rect 3249 14569 3283 14603
rect 7481 14569 7515 14603
rect 11437 14569 11471 14603
rect 12541 14569 12575 14603
rect 12725 14569 12759 14603
rect 14749 14569 14783 14603
rect 5641 14501 5675 14535
rect 10241 14501 10275 14535
rect 1869 14433 1903 14467
rect 4261 14433 4295 14467
rect 9229 14433 9263 14467
rect 10885 14433 10919 14467
rect 13369 14433 13403 14467
rect 4528 14365 4562 14399
rect 6101 14365 6135 14399
rect 8033 14365 8067 14399
rect 8953 14365 8987 14399
rect 10701 14365 10735 14399
rect 11621 14365 11655 14399
rect 11805 14365 11839 14399
rect 11897 14365 11931 14399
rect 13277 14365 13311 14399
rect 13461 14365 13495 14399
rect 14289 14365 14323 14399
rect 14933 14365 14967 14399
rect 15393 14365 15427 14399
rect 15577 14365 15611 14399
rect 2114 14297 2148 14331
rect 6368 14297 6402 14331
rect 8217 14297 8251 14331
rect 12357 14297 12391 14331
rect 10609 14229 10643 14263
rect 12541 14229 12575 14263
rect 14105 14229 14139 14263
rect 15485 14229 15519 14263
rect 5181 14025 5215 14059
rect 10287 14025 10321 14059
rect 12909 14025 12943 14059
rect 1777 13957 1811 13991
rect 1869 13957 1903 13991
rect 7297 13957 7331 13991
rect 14749 13957 14783 13991
rect 15669 13957 15703 13991
rect 2605 13889 2639 13923
rect 4997 13889 5031 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 7113 13889 7147 13923
rect 7389 13889 7423 13923
rect 7849 13889 7883 13923
rect 11529 13889 11563 13923
rect 11713 13889 11747 13923
rect 11989 13889 12023 13923
rect 12541 13889 12575 13923
rect 12725 13889 12759 13923
rect 13001 13889 13035 13923
rect 13553 13889 13587 13923
rect 13737 13889 13771 13923
rect 14381 13889 14415 13923
rect 14565 13889 14599 13923
rect 2053 13821 2087 13855
rect 6929 13821 6963 13855
rect 10057 13821 10091 13855
rect 11897 13821 11931 13855
rect 13921 13821 13955 13855
rect 1409 13753 1443 13787
rect 4353 13753 4387 13787
rect 11805 13753 11839 13787
rect 15853 13753 15887 13787
rect 2868 13685 2902 13719
rect 5641 13685 5675 13719
rect 9137 13685 9171 13719
rect 3249 13481 3283 13515
rect 5549 13481 5583 13515
rect 12081 13481 12115 13515
rect 12909 13481 12943 13515
rect 15669 13481 15703 13515
rect 15025 13413 15059 13447
rect 1777 13345 1811 13379
rect 4077 13345 4111 13379
rect 15761 13345 15795 13379
rect 1501 13277 1535 13311
rect 3801 13277 3835 13311
rect 6009 13277 6043 13311
rect 6193 13277 6227 13311
rect 6653 13277 6687 13311
rect 8401 13277 8435 13311
rect 9321 13277 9355 13311
rect 11529 13277 11563 13311
rect 11713 13277 11747 13311
rect 11897 13277 11931 13311
rect 12541 13277 12575 13311
rect 14289 13277 14323 13311
rect 14565 13277 14599 13311
rect 15209 13277 15243 13311
rect 15669 13277 15703 13311
rect 11069 13209 11103 13243
rect 11805 13209 11839 13243
rect 14105 13209 14139 13243
rect 6101 13141 6135 13175
rect 12909 13141 12943 13175
rect 13093 13141 13127 13175
rect 14473 13141 14507 13175
rect 16037 13141 16071 13175
rect 2237 12937 2271 12971
rect 4813 12937 4847 12971
rect 11529 12937 11563 12971
rect 11989 12937 12023 12971
rect 12725 12937 12759 12971
rect 13093 12937 13127 12971
rect 15485 12937 15519 12971
rect 5457 12869 5491 12903
rect 5549 12869 5583 12903
rect 11897 12869 11931 12903
rect 14289 12869 14323 12903
rect 1777 12801 1811 12835
rect 2053 12801 2087 12835
rect 2513 12801 2547 12835
rect 2973 12801 3007 12835
rect 5273 12801 5307 12835
rect 5641 12801 5675 12835
rect 6377 12801 6411 12835
rect 7849 12801 7883 12835
rect 9413 12801 9447 12835
rect 10149 12801 10183 12835
rect 10793 12801 10827 12835
rect 10977 12801 11011 12835
rect 14105 12801 14139 12835
rect 14381 12801 14415 12835
rect 15301 12801 15335 12835
rect 15577 12801 15611 12835
rect 3157 12733 3191 12767
rect 3893 12733 3927 12767
rect 4031 12733 4065 12767
rect 4169 12733 4203 12767
rect 6653 12733 6687 12767
rect 12081 12733 12115 12767
rect 13185 12733 13219 12767
rect 13277 12733 13311 12767
rect 3617 12665 3651 12699
rect 10793 12665 10827 12699
rect 5825 12597 5859 12631
rect 10241 12597 10275 12631
rect 13921 12597 13955 12631
rect 15117 12597 15151 12631
rect 5641 12393 5675 12427
rect 9045 12393 9079 12427
rect 12909 12325 12943 12359
rect 13369 12325 13403 12359
rect 1409 12257 1443 12291
rect 1593 12257 1627 12291
rect 2053 12257 2087 12291
rect 2467 12257 2501 12291
rect 3985 12257 4019 12291
rect 4445 12257 4479 12291
rect 4721 12257 4755 12291
rect 4997 12257 5031 12291
rect 2329 12189 2363 12223
rect 2605 12189 2639 12223
rect 3801 12189 3835 12223
rect 4838 12189 4872 12223
rect 9229 12189 9263 12223
rect 9689 12189 9723 12223
rect 11529 12189 11563 12223
rect 13553 12189 13587 12223
rect 14289 12189 14323 12223
rect 14565 12189 14599 12223
rect 15209 12189 15243 12223
rect 15485 12189 15519 12223
rect 15945 12189 15979 12223
rect 3249 12121 3283 12155
rect 6653 12121 6687 12155
rect 9956 12121 9990 12155
rect 11796 12121 11830 12155
rect 14105 12121 14139 12155
rect 14473 12121 14507 12155
rect 7941 12053 7975 12087
rect 11069 12053 11103 12087
rect 15025 12053 15059 12087
rect 15393 12053 15427 12087
rect 16129 12053 16163 12087
rect 4721 11849 4755 11883
rect 9689 11849 9723 11883
rect 10609 11849 10643 11883
rect 13921 11849 13955 11883
rect 15393 11849 15427 11883
rect 8401 11781 8435 11815
rect 14749 11781 14783 11815
rect 15761 11781 15795 11815
rect 1593 11713 1627 11747
rect 3065 11713 3099 11747
rect 4077 11713 4111 11747
rect 5181 11713 5215 11747
rect 5457 11713 5491 11747
rect 5641 11713 5675 11747
rect 6561 11713 6595 11747
rect 6828 11713 6862 11747
rect 10793 11713 10827 11747
rect 11785 11713 11819 11747
rect 13369 11713 13403 11747
rect 13553 11713 13587 11747
rect 13645 11713 13679 11747
rect 13737 11713 13771 11747
rect 15577 11713 15611 11747
rect 15853 11713 15887 11747
rect 1869 11645 1903 11679
rect 2881 11645 2915 11679
rect 3801 11645 3835 11679
rect 3939 11645 3973 11679
rect 5825 11645 5859 11679
rect 11529 11645 11563 11679
rect 3525 11577 3559 11611
rect 12909 11577 12943 11611
rect 14381 11577 14415 11611
rect 14933 11577 14967 11611
rect 7941 11509 7975 11543
rect 14771 11509 14805 11543
rect 12173 11305 12207 11339
rect 13553 11305 13587 11339
rect 3249 11237 3283 11271
rect 6193 11237 6227 11271
rect 14657 11237 14691 11271
rect 1501 11169 1535 11203
rect 4445 11169 4479 11203
rect 8953 11169 8987 11203
rect 3801 11101 3835 11135
rect 8401 11101 8435 11135
rect 10793 11101 10827 11135
rect 13001 11101 13035 11135
rect 13185 11101 13219 11135
rect 13277 11101 13311 11135
rect 13393 11101 13427 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 14473 11101 14507 11135
rect 15301 11101 15335 11135
rect 15485 11101 15519 11135
rect 15577 11101 15611 11135
rect 1777 11033 1811 11067
rect 3893 11033 3927 11067
rect 4721 11033 4755 11067
rect 6653 11033 6687 11067
rect 9220 11033 9254 11067
rect 11060 11033 11094 11067
rect 14381 11033 14415 11067
rect 10333 10965 10367 10999
rect 15117 10965 15151 10999
rect 1777 10761 1811 10795
rect 2053 10761 2087 10795
rect 5181 10761 5215 10795
rect 12909 10761 12943 10795
rect 15025 10761 15059 10795
rect 7849 10693 7883 10727
rect 11796 10693 11830 10727
rect 13737 10693 13771 10727
rect 14657 10693 14691 10727
rect 14749 10693 14783 10727
rect 15853 10693 15887 10727
rect 1409 10625 1443 10659
rect 1894 10625 1928 10659
rect 2513 10625 2547 10659
rect 2881 10625 2915 10659
rect 4307 10625 4341 10659
rect 6653 10625 6687 10659
rect 10149 10625 10183 10659
rect 13553 10625 13587 10659
rect 13644 10625 13678 10659
rect 13921 10625 13955 10659
rect 14013 10625 14047 10659
rect 14473 10625 14507 10659
rect 14841 10625 14875 10659
rect 15669 10625 15703 10659
rect 15945 10625 15979 10659
rect 1685 10557 1719 10591
rect 5273 10557 5307 10591
rect 5365 10557 5399 10591
rect 6377 10557 6411 10591
rect 10425 10557 10459 10591
rect 11529 10557 11563 10591
rect 13369 10489 13403 10523
rect 15485 10489 15519 10523
rect 4813 10421 4847 10455
rect 9137 10421 9171 10455
rect 3893 10217 3927 10251
rect 8125 10217 8159 10251
rect 11713 10217 11747 10251
rect 15761 10149 15795 10183
rect 1501 10081 1535 10115
rect 3249 10081 3283 10115
rect 4721 10081 4755 10115
rect 9413 10081 9447 10115
rect 15669 10081 15703 10115
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 4445 10013 4479 10047
rect 6653 10013 6687 10047
rect 9137 10013 9171 10047
rect 12725 10013 12759 10047
rect 13001 10013 13035 10047
rect 14565 10013 14599 10047
rect 14749 10013 14783 10047
rect 14913 10013 14947 10047
rect 15577 10013 15611 10047
rect 15853 10013 15887 10047
rect 1777 9945 1811 9979
rect 10425 9945 10459 9979
rect 14657 9945 14691 9979
rect 15209 9945 15243 9979
rect 6193 9877 6227 9911
rect 14381 9877 14415 9911
rect 15393 9877 15427 9911
rect 14749 9673 14783 9707
rect 9229 9605 9263 9639
rect 2973 9537 3007 9571
rect 3709 9537 3743 9571
rect 4077 9537 4111 9571
rect 5089 9537 5123 9571
rect 6561 9537 6595 9571
rect 7021 9537 7055 9571
rect 11529 9537 11563 9571
rect 11796 9537 11830 9571
rect 13625 9537 13659 9571
rect 15393 9537 15427 9571
rect 15577 9537 15611 9571
rect 15669 9537 15703 9571
rect 2053 9469 2087 9503
rect 2329 9469 2363 9503
rect 2605 9469 2639 9503
rect 3801 9469 3835 9503
rect 3985 9469 4019 9503
rect 5365 9469 5399 9503
rect 13369 9469 13403 9503
rect 2881 9401 2915 9435
rect 5273 9401 5307 9435
rect 8309 9401 8343 9435
rect 12909 9401 12943 9435
rect 5181 9333 5215 9367
rect 6377 9333 6411 9367
rect 10517 9333 10551 9367
rect 15209 9333 15243 9367
rect 3249 9129 3283 9163
rect 6285 9129 6319 9163
rect 8401 9129 8435 9163
rect 14105 9129 14139 9163
rect 1501 8993 1535 9027
rect 7021 8993 7055 9027
rect 11529 8993 11563 9027
rect 14289 8993 14323 9027
rect 14381 8993 14415 9027
rect 14473 8993 14507 9027
rect 3801 8925 3835 8959
rect 3985 8925 4019 8959
rect 4169 8925 4203 8959
rect 4813 8925 4847 8959
rect 9321 8925 9355 8959
rect 13369 8925 13403 8959
rect 13461 8925 13495 8959
rect 14565 8925 14599 8959
rect 15301 8925 15335 8959
rect 15577 8925 15611 8959
rect 1777 8857 1811 8891
rect 4077 8857 4111 8891
rect 7288 8857 7322 8891
rect 11796 8857 11830 8891
rect 15117 8857 15151 8891
rect 15485 8857 15519 8891
rect 4353 8789 4387 8823
rect 10793 8789 10827 8823
rect 12909 8789 12943 8823
rect 3341 8585 3375 8619
rect 13369 8585 13403 8619
rect 15209 8585 15243 8619
rect 13737 8517 13771 8551
rect 3801 8449 3835 8483
rect 8861 8449 8895 8483
rect 10425 8449 10459 8483
rect 11529 8449 11563 8483
rect 11796 8449 11830 8483
rect 14565 8449 14599 8483
rect 15577 8449 15611 8483
rect 15853 8449 15887 8483
rect 1593 8381 1627 8415
rect 1869 8381 1903 8415
rect 4077 8381 4111 8415
rect 5549 8381 5583 8415
rect 6377 8381 6411 8415
rect 6653 8381 6687 8415
rect 13829 8381 13863 8415
rect 14013 8381 14047 8415
rect 14657 8381 14691 8415
rect 15669 8381 15703 8415
rect 14933 8313 14967 8347
rect 3709 8245 3743 8279
rect 8125 8245 8159 8279
rect 12909 8245 12943 8279
rect 15577 8245 15611 8279
rect 16037 8245 16071 8279
rect 15117 8041 15151 8075
rect 6745 7973 6779 8007
rect 1501 7905 1535 7939
rect 1777 7905 1811 7939
rect 9597 7905 9631 7939
rect 14197 7905 14231 7939
rect 3801 7837 3835 7871
rect 4077 7837 4111 7871
rect 7481 7837 7515 7871
rect 7665 7837 7699 7871
rect 7941 7837 7975 7871
rect 12633 7837 12667 7871
rect 12909 7837 12943 7871
rect 14289 7837 14323 7871
rect 15301 7837 15335 7871
rect 15485 7837 15519 7871
rect 15577 7837 15611 7871
rect 5273 7769 5307 7803
rect 10425 7769 10459 7803
rect 3249 7701 3283 7735
rect 7849 7701 7883 7735
rect 8953 7701 8987 7735
rect 9321 7701 9355 7735
rect 9413 7701 9447 7735
rect 11713 7701 11747 7735
rect 14657 7701 14691 7735
rect 4077 7429 4111 7463
rect 5825 7429 5859 7463
rect 7849 7429 7883 7463
rect 12633 7429 12667 7463
rect 1869 7361 1903 7395
rect 7021 7361 7055 7395
rect 7113 7361 7147 7395
rect 10609 7361 10643 7395
rect 10885 7361 10919 7395
rect 11805 7361 11839 7395
rect 12081 7361 12115 7395
rect 15301 7361 15335 7395
rect 15485 7361 15519 7395
rect 15577 7361 15611 7395
rect 2145 7293 2179 7327
rect 7205 7293 7239 7327
rect 10793 7293 10827 7327
rect 11713 7293 11747 7327
rect 12173 7293 12207 7327
rect 15117 7293 15151 7327
rect 10701 7225 10735 7259
rect 11529 7225 11563 7259
rect 3617 7157 3651 7191
rect 6653 7157 6687 7191
rect 9137 7157 9171 7191
rect 10425 7157 10459 7191
rect 13921 7157 13955 7191
rect 1764 6953 1798 6987
rect 11069 6953 11103 6987
rect 9137 6885 9171 6919
rect 12909 6885 12943 6919
rect 15301 6885 15335 6919
rect 1501 6817 1535 6851
rect 6837 6817 6871 6851
rect 9229 6817 9263 6851
rect 9689 6817 9723 6851
rect 3985 6749 4019 6783
rect 4261 6749 4295 6783
rect 5273 6749 5307 6783
rect 8033 6749 8067 6783
rect 8217 6749 8251 6783
rect 8953 6749 8987 6783
rect 9045 6749 9079 6783
rect 9956 6749 9990 6783
rect 11529 6749 11563 6783
rect 11796 6749 11830 6783
rect 13369 6749 13403 6783
rect 14105 6749 14139 6783
rect 14289 6749 14323 6783
rect 14565 6749 14599 6783
rect 15025 6749 15059 6783
rect 15163 6749 15197 6783
rect 15485 6749 15519 6783
rect 16129 6749 16163 6783
rect 8401 6681 8435 6715
rect 15393 6681 15427 6715
rect 3249 6613 3283 6647
rect 13461 6613 13495 6647
rect 14473 6613 14507 6647
rect 15945 6613 15979 6647
rect 5549 6409 5583 6443
rect 6929 6409 6963 6443
rect 8769 6409 8803 6443
rect 14749 6409 14783 6443
rect 14289 6341 14323 6375
rect 1593 6273 1627 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 6653 6273 6687 6307
rect 6745 6273 6779 6307
rect 7389 6273 7423 6307
rect 7656 6273 7690 6307
rect 9229 6273 9263 6307
rect 9496 6273 9530 6307
rect 11785 6273 11819 6307
rect 13553 6273 13587 6307
rect 13737 6273 13771 6307
rect 13829 6273 13863 6307
rect 15209 6273 15243 6307
rect 15393 6273 15427 6307
rect 1869 6205 1903 6239
rect 3801 6205 3835 6239
rect 4077 6205 4111 6239
rect 11529 6205 11563 6239
rect 13369 6137 13403 6171
rect 14565 6137 14599 6171
rect 3341 6069 3375 6103
rect 10609 6069 10643 6103
rect 12909 6069 12943 6103
rect 15209 6069 15243 6103
rect 15577 6069 15611 6103
rect 6745 5865 6779 5899
rect 9321 5865 9355 5899
rect 14105 5865 14139 5899
rect 14473 5865 14507 5899
rect 15853 5865 15887 5899
rect 1501 5729 1535 5763
rect 1777 5729 1811 5763
rect 3985 5729 4019 5763
rect 13001 5729 13035 5763
rect 14197 5729 14231 5763
rect 4261 5661 4295 5695
rect 5273 5661 5307 5695
rect 8033 5661 8067 5695
rect 8217 5661 8251 5695
rect 8309 5661 8343 5695
rect 9505 5661 9539 5695
rect 9827 5661 9861 5695
rect 9965 5661 9999 5695
rect 10258 5661 10292 5695
rect 14105 5661 14139 5695
rect 15301 5661 15335 5695
rect 15853 5661 15887 5695
rect 15945 5661 15979 5695
rect 9594 5593 9628 5627
rect 9689 5593 9723 5627
rect 12633 5593 12667 5627
rect 12817 5593 12851 5627
rect 14933 5593 14967 5627
rect 15117 5593 15151 5627
rect 3249 5525 3283 5559
rect 7849 5525 7883 5559
rect 11529 5525 11563 5559
rect 12265 5525 12299 5559
rect 9229 5321 9263 5355
rect 11529 5321 11563 5355
rect 7941 5253 7975 5287
rect 11897 5253 11931 5287
rect 12817 5253 12851 5287
rect 15361 5253 15395 5287
rect 15577 5253 15611 5287
rect 1409 5185 1443 5219
rect 1685 5185 1719 5219
rect 2237 5185 2271 5219
rect 2493 5185 2527 5219
rect 4077 5185 4111 5219
rect 6377 5185 6411 5219
rect 6565 5191 6599 5225
rect 6884 5185 6918 5219
rect 10333 5185 10367 5219
rect 10609 5185 10643 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 14565 5185 14599 5219
rect 1777 5117 1811 5151
rect 6653 5117 6687 5151
rect 6745 5117 6779 5151
rect 7113 5117 7147 5151
rect 10149 5117 10183 5151
rect 10425 5117 10459 5151
rect 10517 5049 10551 5083
rect 14841 5049 14875 5083
rect 3617 4981 3651 5015
rect 5365 4981 5399 5015
rect 15209 4981 15243 5015
rect 15393 4981 15427 5015
rect 12633 4777 12667 4811
rect 13001 4777 13035 4811
rect 14289 4777 14323 4811
rect 15853 4777 15887 4811
rect 15945 4777 15979 4811
rect 2605 4709 2639 4743
rect 8309 4709 8343 4743
rect 8953 4709 8987 4743
rect 15025 4709 15059 4743
rect 1501 4641 1535 4675
rect 7941 4641 7975 4675
rect 9413 4641 9447 4675
rect 12725 4641 12759 4675
rect 16037 4641 16071 4675
rect 1593 4573 1627 4607
rect 2421 4573 2455 4607
rect 2697 4573 2731 4607
rect 2973 4573 3007 4607
rect 3157 4573 3191 4607
rect 3801 4573 3835 4607
rect 4077 4573 4111 4607
rect 5273 4573 5307 4607
rect 7021 4573 7055 4607
rect 9137 4573 9171 4607
rect 9229 4573 9263 4607
rect 9321 4573 9355 4607
rect 10425 4573 10459 4607
rect 12633 4573 12667 4607
rect 14933 4573 14967 4607
rect 15117 4573 15151 4607
rect 15761 4573 15795 4607
rect 12173 4505 12207 4539
rect 14105 4505 14139 4539
rect 14321 4505 14355 4539
rect 1961 4437 1995 4471
rect 8401 4437 8435 4471
rect 14473 4437 14507 4471
rect 11897 4233 11931 4267
rect 1777 4165 1811 4199
rect 2872 4165 2906 4199
rect 1409 4097 1443 4131
rect 4445 4097 4479 4131
rect 4701 4097 4735 4131
rect 6561 4097 6595 4131
rect 7113 4097 7147 4131
rect 7380 4097 7414 4131
rect 9229 4097 9263 4131
rect 11713 4097 11747 4131
rect 11989 4097 12023 4131
rect 13093 4097 13127 4131
rect 13185 4097 13219 4131
rect 13829 4097 13863 4131
rect 14105 4097 14139 4131
rect 14749 4097 14783 4131
rect 15853 4097 15887 4131
rect 16037 4097 16071 4131
rect 16129 4097 16163 4131
rect 2605 4029 2639 4063
rect 10793 4029 10827 4063
rect 11529 4029 11563 4063
rect 13369 4029 13403 4063
rect 14933 4029 14967 4063
rect 3985 3961 4019 3995
rect 5825 3961 5859 3995
rect 6377 3961 6411 3995
rect 13921 3961 13955 3995
rect 1777 3893 1811 3927
rect 1961 3893 1995 3927
rect 8493 3893 8527 3927
rect 15853 3893 15887 3927
rect 6745 3689 6779 3723
rect 10977 3689 11011 3723
rect 13185 3689 13219 3723
rect 14289 3689 14323 3723
rect 2973 3621 3007 3655
rect 8033 3621 8067 3655
rect 11713 3621 11747 3655
rect 15485 3621 15519 3655
rect 1685 3553 1719 3587
rect 1961 3553 1995 3587
rect 4077 3553 4111 3587
rect 8953 3553 8987 3587
rect 14933 3553 14967 3587
rect 3157 3485 3191 3519
rect 3249 3485 3283 3519
rect 3801 3485 3835 3519
rect 5273 3485 5307 3519
rect 7481 3485 7515 3519
rect 7665 3485 7699 3519
rect 7849 3485 7883 3519
rect 9209 3485 9243 3519
rect 11621 3485 11655 3519
rect 11897 3485 11931 3519
rect 12449 3485 12483 3519
rect 12725 3485 12759 3519
rect 13369 3485 13403 3519
rect 14841 3485 14875 3519
rect 15669 3485 15703 3519
rect 2973 3417 3007 3451
rect 7757 3417 7791 3451
rect 10793 3417 10827 3451
rect 10993 3417 11027 3451
rect 14197 3417 14231 3451
rect 10333 3349 10367 3383
rect 11161 3349 11195 3383
rect 12547 3349 12581 3383
rect 12633 3349 12667 3383
rect 1593 3145 1627 3179
rect 10241 3145 10275 3179
rect 11897 3145 11931 3179
rect 13369 3145 13403 3179
rect 15301 3145 15335 3179
rect 4712 3077 4746 3111
rect 6745 3077 6779 3111
rect 9597 3077 9631 3111
rect 10057 3077 10091 3111
rect 11529 3077 11563 3111
rect 11713 3077 11747 3111
rect 13921 3077 13955 3111
rect 14105 3077 14139 3111
rect 1961 3009 1995 3043
rect 2605 3009 2639 3043
rect 2872 3009 2906 3043
rect 4445 3009 4479 3043
rect 6377 3009 6411 3043
rect 6525 3009 6559 3043
rect 6653 3009 6687 3043
rect 6883 3009 6917 3043
rect 7849 3009 7883 3043
rect 12357 3009 12391 3043
rect 12633 3009 12667 3043
rect 13185 3009 13219 3043
rect 13461 3009 13495 3043
rect 14197 3009 14231 3043
rect 14657 3009 14691 3043
rect 14841 3009 14875 3043
rect 15485 3009 15519 3043
rect 15945 3009 15979 3043
rect 1777 2941 1811 2975
rect 1869 2941 1903 2975
rect 2053 2941 2087 2975
rect 3985 2873 4019 2907
rect 5825 2873 5859 2907
rect 12449 2873 12483 2907
rect 13185 2873 13219 2907
rect 16129 2873 16163 2907
rect 7021 2805 7055 2839
rect 10241 2805 10275 2839
rect 10425 2805 10459 2839
rect 13921 2805 13955 2839
rect 14657 2805 14691 2839
rect 7573 2601 7607 2635
rect 8033 2601 8067 2635
rect 11713 2601 11747 2635
rect 14289 2601 14323 2635
rect 15853 2601 15887 2635
rect 3801 2533 3835 2567
rect 11161 2533 11195 2567
rect 13369 2533 13403 2567
rect 1409 2465 1443 2499
rect 1685 2465 1719 2499
rect 2789 2465 2823 2499
rect 4445 2465 4479 2499
rect 7021 2465 7055 2499
rect 12817 2465 12851 2499
rect 2881 2397 2915 2431
rect 7481 2397 7515 2431
rect 7757 2397 7791 2431
rect 9137 2397 9171 2431
rect 9413 2397 9447 2431
rect 10057 2397 10091 2431
rect 10333 2397 10367 2431
rect 10793 2397 10827 2431
rect 10977 2397 11011 2431
rect 11621 2397 11655 2431
rect 11805 2397 11839 2431
rect 12541 2397 12575 2431
rect 12725 2397 12759 2431
rect 13277 2397 13311 2431
rect 13553 2397 13587 2431
rect 14197 2397 14231 2431
rect 15025 2397 15059 2431
rect 15853 2397 15887 2431
rect 16037 2397 16071 2431
rect 4261 2329 4295 2363
rect 5273 2329 5307 2363
rect 13461 2329 13495 2363
rect 3249 2261 3283 2295
rect 4169 2261 4203 2295
rect 8953 2261 8987 2295
rect 9321 2261 9355 2295
rect 9873 2261 9907 2295
rect 10241 2261 10275 2295
rect 14841 2261 14875 2295
rect 3065 2057 3099 2091
rect 3801 2057 3835 2091
rect 5825 2057 5859 2091
rect 12725 2057 12759 2091
rect 14933 2057 14967 2091
rect 15577 2057 15611 2091
rect 4169 1989 4203 2023
rect 5457 1989 5491 2023
rect 6377 1989 6411 2023
rect 10241 1989 10275 2023
rect 10885 1989 10919 2023
rect 14013 1989 14047 2023
rect 14229 1989 14263 2023
rect 2053 1921 2087 1955
rect 4261 1921 4295 1955
rect 5273 1921 5307 1955
rect 5549 1921 5583 1955
rect 5641 1921 5675 1955
rect 6561 1921 6595 1955
rect 6653 1921 6687 1955
rect 7113 1921 7147 1955
rect 7380 1921 7414 1955
rect 8953 1921 8987 1955
rect 9873 1921 9907 1955
rect 10057 1921 10091 1955
rect 10333 1921 10367 1955
rect 10793 1921 10827 1955
rect 10977 1921 11011 1955
rect 11529 1921 11563 1955
rect 11713 1921 11747 1955
rect 11897 1921 11931 1955
rect 12357 1921 12391 1955
rect 12449 1921 12483 1955
rect 13185 1921 13219 1955
rect 13369 1921 13403 1955
rect 14841 1921 14875 1955
rect 15025 1921 15059 1955
rect 15485 1921 15519 1955
rect 1869 1853 1903 1887
rect 1961 1853 1995 1887
rect 2145 1853 2179 1887
rect 2697 1853 2731 1887
rect 4445 1853 4479 1887
rect 3249 1785 3283 1819
rect 8493 1785 8527 1819
rect 13277 1785 13311 1819
rect 1685 1717 1719 1751
rect 3065 1717 3099 1751
rect 6653 1717 6687 1751
rect 9229 1717 9263 1751
rect 9413 1717 9447 1751
rect 12541 1717 12575 1751
rect 14197 1717 14231 1751
rect 14381 1717 14415 1751
rect 1869 1513 1903 1547
rect 2789 1513 2823 1547
rect 4169 1513 4203 1547
rect 6561 1513 6595 1547
rect 8217 1513 8251 1547
rect 8953 1513 8987 1547
rect 10057 1513 10091 1547
rect 11713 1513 11747 1547
rect 13277 1513 13311 1547
rect 14289 1513 14323 1547
rect 14473 1513 14507 1547
rect 4905 1445 4939 1479
rect 4997 1445 5031 1479
rect 5641 1445 5675 1479
rect 7665 1445 7699 1479
rect 12449 1445 12483 1479
rect 15209 1445 15243 1479
rect 3801 1377 3835 1411
rect 2053 1309 2087 1343
rect 2237 1309 2271 1343
rect 2329 1309 2363 1343
rect 2973 1309 3007 1343
rect 3249 1309 3283 1343
rect 3985 1309 4019 1343
rect 4813 1309 4847 1343
rect 5089 1309 5123 1343
rect 5825 1309 5859 1343
rect 6837 1309 6871 1343
rect 8401 1309 8435 1343
rect 9137 1309 9171 1343
rect 9413 1309 9447 1343
rect 10793 1309 10827 1343
rect 12357 1309 12391 1343
rect 12633 1309 12667 1343
rect 13185 1309 13219 1343
rect 13461 1309 13495 1343
rect 15025 1309 15059 1343
rect 15853 1309 15887 1343
rect 6377 1241 6411 1275
rect 6561 1241 6595 1275
rect 7297 1241 7331 1275
rect 9321 1241 9355 1275
rect 9873 1241 9907 1275
rect 10089 1241 10123 1275
rect 11529 1241 11563 1275
rect 14105 1241 14139 1275
rect 3157 1173 3191 1207
rect 4629 1173 4663 1207
rect 7757 1173 7791 1207
rect 10241 1173 10275 1207
rect 10885 1173 10919 1207
rect 11729 1173 11763 1207
rect 11897 1173 11931 1207
rect 14305 1173 14339 1207
rect 15669 1173 15703 1207
<< metal1 >>
rect 1104 22874 16836 22896
rect 1104 22822 4898 22874
rect 4950 22822 4962 22874
rect 5014 22822 5026 22874
rect 5078 22822 5090 22874
rect 5142 22822 5154 22874
rect 5206 22822 8846 22874
rect 8898 22822 8910 22874
rect 8962 22822 8974 22874
rect 9026 22822 9038 22874
rect 9090 22822 9102 22874
rect 9154 22822 12794 22874
rect 12846 22822 12858 22874
rect 12910 22822 12922 22874
rect 12974 22822 12986 22874
rect 13038 22822 13050 22874
rect 13102 22822 16836 22874
rect 1104 22800 16836 22822
rect 1397 22627 1455 22633
rect 1397 22593 1409 22627
rect 1443 22593 1455 22627
rect 1397 22587 1455 22593
rect 1581 22627 1639 22633
rect 1581 22593 1593 22627
rect 1627 22624 1639 22627
rect 14182 22624 14188 22636
rect 1627 22596 14188 22624
rect 1627 22593 1639 22596
rect 1581 22587 1639 22593
rect 1412 22556 1440 22587
rect 14182 22584 14188 22596
rect 14240 22584 14246 22636
rect 1412 22528 1992 22556
rect 1486 22488 1492 22500
rect 1447 22460 1492 22488
rect 1486 22448 1492 22460
rect 1544 22448 1550 22500
rect 1964 22429 1992 22528
rect 1949 22423 2007 22429
rect 1949 22389 1961 22423
rect 1995 22420 2007 22423
rect 16942 22420 16948 22432
rect 1995 22392 16948 22420
rect 1995 22389 2007 22392
rect 1949 22383 2007 22389
rect 16942 22380 16948 22392
rect 17000 22380 17006 22432
rect 1104 22330 16836 22352
rect 1104 22278 2924 22330
rect 2976 22278 2988 22330
rect 3040 22278 3052 22330
rect 3104 22278 3116 22330
rect 3168 22278 3180 22330
rect 3232 22278 6872 22330
rect 6924 22278 6936 22330
rect 6988 22278 7000 22330
rect 7052 22278 7064 22330
rect 7116 22278 7128 22330
rect 7180 22278 10820 22330
rect 10872 22278 10884 22330
rect 10936 22278 10948 22330
rect 11000 22278 11012 22330
rect 11064 22278 11076 22330
rect 11128 22278 14768 22330
rect 14820 22278 14832 22330
rect 14884 22278 14896 22330
rect 14948 22278 14960 22330
rect 15012 22278 15024 22330
rect 15076 22278 16836 22330
rect 1104 22256 16836 22278
rect 1578 22216 1584 22228
rect 1539 22188 1584 22216
rect 1578 22176 1584 22188
rect 1636 22176 1642 22228
rect 2774 22148 2780 22160
rect 2735 22120 2780 22148
rect 2774 22108 2780 22120
rect 2832 22108 2838 22160
rect 8018 22080 8024 22092
rect 2746 22052 8024 22080
rect 1397 22015 1455 22021
rect 1397 21981 1409 22015
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 2317 22015 2375 22021
rect 2317 21981 2329 22015
rect 2363 22012 2375 22015
rect 2746 22012 2774 22052
rect 8018 22040 8024 22052
rect 8076 22040 8082 22092
rect 2363 21984 2774 22012
rect 2961 22015 3019 22021
rect 2363 21981 2375 21984
rect 2317 21975 2375 21981
rect 2961 21981 2973 22015
rect 3007 22012 3019 22015
rect 3878 22012 3884 22024
rect 3007 21984 3884 22012
rect 3007 21981 3019 21984
rect 2961 21975 3019 21981
rect 1412 21944 1440 21975
rect 3878 21972 3884 21984
rect 3936 21972 3942 22024
rect 8570 21944 8576 21956
rect 1412 21916 8576 21944
rect 8570 21904 8576 21916
rect 8628 21904 8634 21956
rect 2133 21879 2191 21885
rect 2133 21845 2145 21879
rect 2179 21876 2191 21879
rect 6730 21876 6736 21888
rect 2179 21848 6736 21876
rect 2179 21845 2191 21848
rect 2133 21839 2191 21845
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 1104 21786 16836 21808
rect 1104 21734 4898 21786
rect 4950 21734 4962 21786
rect 5014 21734 5026 21786
rect 5078 21734 5090 21786
rect 5142 21734 5154 21786
rect 5206 21734 8846 21786
rect 8898 21734 8910 21786
rect 8962 21734 8974 21786
rect 9026 21734 9038 21786
rect 9090 21734 9102 21786
rect 9154 21734 12794 21786
rect 12846 21734 12858 21786
rect 12910 21734 12922 21786
rect 12974 21734 12986 21786
rect 13038 21734 13050 21786
rect 13102 21734 16836 21786
rect 1104 21712 16836 21734
rect 382 21632 388 21684
rect 440 21672 446 21684
rect 440 21644 3832 21672
rect 440 21632 446 21644
rect 1504 21576 3096 21604
rect 1504 21545 1532 21576
rect 1489 21539 1547 21545
rect 1489 21505 1501 21539
rect 1535 21505 1547 21539
rect 1489 21499 1547 21505
rect 2225 21539 2283 21545
rect 2225 21505 2237 21539
rect 2271 21536 2283 21539
rect 2271 21508 2774 21536
rect 2271 21505 2283 21508
rect 2225 21499 2283 21505
rect 2746 21400 2774 21508
rect 2961 21403 3019 21409
rect 2961 21400 2973 21403
rect 2746 21372 2973 21400
rect 2961 21369 2973 21372
rect 3007 21369 3019 21403
rect 3068 21400 3096 21576
rect 3804 21545 3832 21644
rect 3145 21539 3203 21545
rect 3145 21505 3157 21539
rect 3191 21505 3203 21539
rect 3145 21499 3203 21505
rect 3789 21539 3847 21545
rect 3789 21505 3801 21539
rect 3835 21505 3847 21539
rect 3789 21499 3847 21505
rect 3160 21468 3188 21499
rect 4062 21468 4068 21480
rect 3160 21440 4068 21468
rect 4062 21428 4068 21440
rect 4120 21428 4126 21480
rect 9306 21400 9312 21412
rect 3068 21372 9312 21400
rect 2961 21363 3019 21369
rect 9306 21360 9312 21372
rect 9364 21360 9370 21412
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 1673 21335 1731 21341
rect 1673 21332 1685 21335
rect 1452 21304 1685 21332
rect 1452 21292 1458 21304
rect 1673 21301 1685 21304
rect 1719 21301 1731 21335
rect 1673 21295 1731 21301
rect 2409 21335 2467 21341
rect 2409 21301 2421 21335
rect 2455 21332 2467 21335
rect 3418 21332 3424 21344
rect 2455 21304 3424 21332
rect 2455 21301 2467 21304
rect 2409 21295 2467 21301
rect 3418 21292 3424 21304
rect 3476 21292 3482 21344
rect 3602 21332 3608 21344
rect 3563 21304 3608 21332
rect 3602 21292 3608 21304
rect 3660 21292 3666 21344
rect 1104 21242 16836 21264
rect 1104 21190 2924 21242
rect 2976 21190 2988 21242
rect 3040 21190 3052 21242
rect 3104 21190 3116 21242
rect 3168 21190 3180 21242
rect 3232 21190 6872 21242
rect 6924 21190 6936 21242
rect 6988 21190 7000 21242
rect 7052 21190 7064 21242
rect 7116 21190 7128 21242
rect 7180 21190 10820 21242
rect 10872 21190 10884 21242
rect 10936 21190 10948 21242
rect 11000 21190 11012 21242
rect 11064 21190 11076 21242
rect 11128 21190 14768 21242
rect 14820 21190 14832 21242
rect 14884 21190 14896 21242
rect 14948 21190 14960 21242
rect 15012 21190 15024 21242
rect 15076 21190 16836 21242
rect 1104 21168 16836 21190
rect 2406 21128 2412 21140
rect 2367 21100 2412 21128
rect 2406 21088 2412 21100
rect 2464 21088 2470 21140
rect 1486 20924 1492 20936
rect 1447 20896 1492 20924
rect 1486 20884 1492 20896
rect 1544 20884 1550 20936
rect 2222 20924 2228 20936
rect 2183 20896 2228 20924
rect 2222 20884 2228 20896
rect 2280 20884 2286 20936
rect 2774 20884 2780 20936
rect 2832 20924 2838 20936
rect 2961 20927 3019 20933
rect 2961 20924 2973 20927
rect 2832 20896 2973 20924
rect 2832 20884 2838 20896
rect 2961 20893 2973 20896
rect 3007 20893 3019 20927
rect 3970 20924 3976 20936
rect 3931 20896 3976 20924
rect 2961 20887 3019 20893
rect 3970 20884 3976 20896
rect 4028 20884 4034 20936
rect 4617 20927 4675 20933
rect 4617 20893 4629 20927
rect 4663 20924 4675 20927
rect 10410 20924 10416 20936
rect 4663 20896 10416 20924
rect 4663 20893 4675 20896
rect 4617 20887 4675 20893
rect 10410 20884 10416 20896
rect 10468 20884 10474 20936
rect 2682 20816 2688 20868
rect 2740 20856 2746 20868
rect 3602 20856 3608 20868
rect 2740 20828 3608 20856
rect 2740 20816 2746 20828
rect 3602 20816 3608 20828
rect 3660 20816 3666 20868
rect 1578 20748 1584 20800
rect 1636 20788 1642 20800
rect 1673 20791 1731 20797
rect 1673 20788 1685 20791
rect 1636 20760 1685 20788
rect 1636 20748 1642 20760
rect 1673 20757 1685 20760
rect 1719 20757 1731 20791
rect 1673 20751 1731 20757
rect 3145 20791 3203 20797
rect 3145 20757 3157 20791
rect 3191 20788 3203 20791
rect 3694 20788 3700 20800
rect 3191 20760 3700 20788
rect 3191 20757 3203 20760
rect 3145 20751 3203 20757
rect 3694 20748 3700 20760
rect 3752 20748 3758 20800
rect 3786 20748 3792 20800
rect 3844 20788 3850 20800
rect 3844 20760 3889 20788
rect 3844 20748 3850 20760
rect 4154 20748 4160 20800
rect 4212 20788 4218 20800
rect 4433 20791 4491 20797
rect 4433 20788 4445 20791
rect 4212 20760 4445 20788
rect 4212 20748 4218 20760
rect 4433 20757 4445 20760
rect 4479 20757 4491 20791
rect 4433 20751 4491 20757
rect 1104 20698 16836 20720
rect 1104 20646 4898 20698
rect 4950 20646 4962 20698
rect 5014 20646 5026 20698
rect 5078 20646 5090 20698
rect 5142 20646 5154 20698
rect 5206 20646 8846 20698
rect 8898 20646 8910 20698
rect 8962 20646 8974 20698
rect 9026 20646 9038 20698
rect 9090 20646 9102 20698
rect 9154 20646 12794 20698
rect 12846 20646 12858 20698
rect 12910 20646 12922 20698
rect 12974 20646 12986 20698
rect 13038 20646 13050 20698
rect 13102 20646 16836 20698
rect 1104 20624 16836 20646
rect 2774 20544 2780 20596
rect 2832 20584 2838 20596
rect 3697 20587 3755 20593
rect 3697 20584 3709 20587
rect 2832 20556 3709 20584
rect 2832 20544 2838 20556
rect 3697 20553 3709 20556
rect 3743 20553 3755 20587
rect 3697 20547 3755 20553
rect 4065 20587 4123 20593
rect 4065 20553 4077 20587
rect 4111 20553 4123 20587
rect 4065 20547 4123 20553
rect 4080 20516 4108 20547
rect 4614 20544 4620 20596
rect 4672 20584 4678 20596
rect 4893 20587 4951 20593
rect 4893 20584 4905 20587
rect 4672 20556 4905 20584
rect 4672 20544 4678 20556
rect 4893 20553 4905 20556
rect 4939 20553 4951 20587
rect 4893 20547 4951 20553
rect 15286 20516 15292 20528
rect 2056 20488 4108 20516
rect 5000 20488 15292 20516
rect 1026 20408 1032 20460
rect 1084 20448 1090 20460
rect 2056 20457 2084 20488
rect 1581 20451 1639 20457
rect 1581 20448 1593 20451
rect 1084 20420 1593 20448
rect 1084 20408 1090 20420
rect 1581 20417 1593 20420
rect 1627 20417 1639 20451
rect 1581 20411 1639 20417
rect 2041 20451 2099 20457
rect 2041 20417 2053 20451
rect 2087 20417 2099 20451
rect 2041 20411 2099 20417
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20448 2835 20451
rect 3142 20448 3148 20460
rect 2823 20420 3148 20448
rect 2823 20417 2835 20420
rect 2777 20411 2835 20417
rect 3142 20408 3148 20420
rect 3200 20408 3206 20460
rect 3513 20451 3571 20457
rect 3513 20417 3525 20451
rect 3559 20448 3571 20451
rect 4154 20448 4160 20460
rect 3559 20420 4160 20448
rect 3559 20417 3571 20420
rect 3513 20411 3571 20417
rect 4154 20408 4160 20420
rect 4212 20408 4218 20460
rect 4246 20408 4252 20460
rect 4304 20448 4310 20460
rect 5000 20448 5028 20488
rect 15286 20476 15292 20488
rect 15344 20476 15350 20528
rect 4304 20420 4349 20448
rect 4540 20420 5028 20448
rect 5077 20451 5135 20457
rect 4304 20408 4310 20420
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20380 3111 20383
rect 3326 20380 3332 20392
rect 3099 20352 3332 20380
rect 3099 20349 3111 20352
rect 3053 20343 3111 20349
rect 3326 20340 3332 20352
rect 3384 20380 3390 20392
rect 4540 20380 4568 20420
rect 5077 20417 5089 20451
rect 5123 20417 5135 20451
rect 5077 20411 5135 20417
rect 5721 20451 5779 20457
rect 5721 20417 5733 20451
rect 5767 20448 5779 20451
rect 9674 20448 9680 20460
rect 5767 20420 9680 20448
rect 5767 20417 5779 20420
rect 5721 20411 5779 20417
rect 3384 20352 4568 20380
rect 4617 20383 4675 20389
rect 3384 20340 3390 20352
rect 4617 20349 4629 20383
rect 4663 20380 4675 20383
rect 5092 20380 5120 20411
rect 9674 20408 9680 20420
rect 9732 20408 9738 20460
rect 17310 20448 17316 20460
rect 12406 20420 17316 20448
rect 12406 20380 12434 20420
rect 17310 20408 17316 20420
rect 17368 20408 17374 20460
rect 4663 20352 12434 20380
rect 4663 20349 4675 20352
rect 4617 20343 4675 20349
rect 2406 20272 2412 20324
rect 2464 20312 2470 20324
rect 2777 20315 2835 20321
rect 2777 20312 2789 20315
rect 2464 20284 2789 20312
rect 2464 20272 2470 20284
rect 2777 20281 2789 20284
rect 2823 20281 2835 20315
rect 2777 20275 2835 20281
rect 2869 20315 2927 20321
rect 2869 20281 2881 20315
rect 2915 20312 2927 20315
rect 3510 20312 3516 20324
rect 2915 20284 3516 20312
rect 2915 20281 2927 20284
rect 2869 20275 2927 20281
rect 3510 20272 3516 20284
rect 3568 20272 3574 20324
rect 4154 20272 4160 20324
rect 4212 20312 4218 20324
rect 16022 20312 16028 20324
rect 4212 20284 16028 20312
rect 4212 20272 4218 20284
rect 16022 20272 16028 20284
rect 16080 20272 16086 20324
rect 1397 20247 1455 20253
rect 1397 20213 1409 20247
rect 1443 20244 1455 20247
rect 1762 20244 1768 20256
rect 1443 20216 1768 20244
rect 1443 20213 1455 20216
rect 1397 20207 1455 20213
rect 1762 20204 1768 20216
rect 1820 20204 1826 20256
rect 1854 20204 1860 20256
rect 1912 20244 1918 20256
rect 2225 20247 2283 20253
rect 2225 20244 2237 20247
rect 1912 20216 2237 20244
rect 1912 20204 1918 20216
rect 2225 20213 2237 20216
rect 2271 20213 2283 20247
rect 2225 20207 2283 20213
rect 2314 20204 2320 20256
rect 2372 20244 2378 20256
rect 4798 20244 4804 20256
rect 2372 20216 4804 20244
rect 2372 20204 2378 20216
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 5537 20247 5595 20253
rect 5537 20213 5549 20247
rect 5583 20244 5595 20247
rect 5718 20244 5724 20256
rect 5583 20216 5724 20244
rect 5583 20213 5595 20216
rect 5537 20207 5595 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 5810 20204 5816 20256
rect 5868 20244 5874 20256
rect 17402 20244 17408 20256
rect 5868 20216 17408 20244
rect 5868 20204 5874 20216
rect 17402 20204 17408 20216
rect 17460 20204 17466 20256
rect 1104 20154 16836 20176
rect 1104 20102 2924 20154
rect 2976 20102 2988 20154
rect 3040 20102 3052 20154
rect 3104 20102 3116 20154
rect 3168 20102 3180 20154
rect 3232 20102 6872 20154
rect 6924 20102 6936 20154
rect 6988 20102 7000 20154
rect 7052 20102 7064 20154
rect 7116 20102 7128 20154
rect 7180 20102 10820 20154
rect 10872 20102 10884 20154
rect 10936 20102 10948 20154
rect 11000 20102 11012 20154
rect 11064 20102 11076 20154
rect 11128 20102 14768 20154
rect 14820 20102 14832 20154
rect 14884 20102 14896 20154
rect 14948 20102 14960 20154
rect 15012 20102 15024 20154
rect 15076 20102 16836 20154
rect 1104 20080 16836 20102
rect 2409 20043 2467 20049
rect 2409 20009 2421 20043
rect 2455 20040 2467 20043
rect 3970 20040 3976 20052
rect 2455 20012 3976 20040
rect 2455 20009 2467 20012
rect 2409 20003 2467 20009
rect 3970 20000 3976 20012
rect 4028 20000 4034 20052
rect 4798 20000 4804 20052
rect 4856 20040 4862 20052
rect 17218 20040 17224 20052
rect 4856 20012 17224 20040
rect 4856 20000 4862 20012
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 3053 19975 3111 19981
rect 3053 19941 3065 19975
rect 3099 19972 3111 19975
rect 3510 19972 3516 19984
rect 3099 19944 3516 19972
rect 3099 19941 3111 19944
rect 3053 19935 3111 19941
rect 3510 19932 3516 19944
rect 3568 19932 3574 19984
rect 3786 19972 3792 19984
rect 3747 19944 3792 19972
rect 3786 19932 3792 19944
rect 3844 19932 3850 19984
rect 5350 19972 5356 19984
rect 5311 19944 5356 19972
rect 5350 19932 5356 19944
rect 5408 19932 5414 19984
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19904 1823 19907
rect 3602 19904 3608 19916
rect 1811 19876 3608 19904
rect 1811 19873 1823 19876
rect 1765 19867 1823 19873
rect 2240 19845 2268 19876
rect 3602 19864 3608 19876
rect 3660 19864 3666 19916
rect 4154 19904 4160 19916
rect 3988 19876 4160 19904
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19805 2191 19839
rect 2133 19799 2191 19805
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19805 2283 19839
rect 2225 19799 2283 19805
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19805 3019 19839
rect 2961 19799 3019 19805
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19836 3295 19839
rect 3326 19836 3332 19848
rect 3283 19808 3332 19836
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 2148 19768 2176 19799
rect 2866 19768 2872 19780
rect 2148 19740 2872 19768
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 2976 19768 3004 19799
rect 3326 19796 3332 19808
rect 3384 19796 3390 19848
rect 3988 19845 4016 19876
rect 4154 19864 4160 19876
rect 4212 19864 4218 19916
rect 6454 19904 6460 19916
rect 5460 19876 6460 19904
rect 3973 19839 4031 19845
rect 3973 19836 3985 19839
rect 3436 19808 3985 19836
rect 3436 19768 3464 19808
rect 3973 19805 3985 19808
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19836 4123 19839
rect 4338 19836 4344 19848
rect 4111 19808 4344 19836
rect 4111 19805 4123 19808
rect 4065 19799 4123 19805
rect 4338 19796 4344 19808
rect 4396 19796 4402 19848
rect 4522 19796 4528 19848
rect 4580 19836 4586 19848
rect 5169 19839 5227 19845
rect 4580 19808 4625 19836
rect 4580 19796 4586 19808
rect 5169 19805 5181 19839
rect 5215 19836 5227 19839
rect 5215 19832 5304 19836
rect 5460 19832 5488 19876
rect 6454 19864 6460 19876
rect 6512 19864 6518 19916
rect 5810 19836 5816 19848
rect 5215 19808 5488 19832
rect 5771 19808 5816 19836
rect 5215 19805 5227 19808
rect 5169 19799 5227 19805
rect 5276 19804 5488 19808
rect 5810 19796 5816 19808
rect 5868 19796 5874 19848
rect 6009 19839 6067 19845
rect 6009 19805 6021 19839
rect 6055 19836 6067 19839
rect 6641 19839 6699 19845
rect 6055 19808 6132 19836
rect 6055 19805 6067 19808
rect 6009 19799 6067 19805
rect 2976 19740 3464 19768
rect 3510 19728 3516 19780
rect 3568 19768 3574 19780
rect 3789 19771 3847 19777
rect 3789 19768 3801 19771
rect 3568 19740 3801 19768
rect 3568 19728 3574 19740
rect 3789 19737 3801 19740
rect 3835 19768 3847 19771
rect 4356 19768 4384 19796
rect 3835 19740 4016 19768
rect 4356 19740 5136 19768
rect 3835 19737 3847 19740
rect 3789 19731 3847 19737
rect 3988 19712 4016 19740
rect 2961 19703 3019 19709
rect 2961 19669 2973 19703
rect 3007 19700 3019 19703
rect 3602 19700 3608 19712
rect 3007 19672 3608 19700
rect 3007 19669 3019 19672
rect 2961 19663 3019 19669
rect 3602 19660 3608 19672
rect 3660 19660 3666 19712
rect 3970 19660 3976 19712
rect 4028 19660 4034 19712
rect 4338 19660 4344 19712
rect 4396 19700 4402 19712
rect 4617 19703 4675 19709
rect 4617 19700 4629 19703
rect 4396 19672 4629 19700
rect 4396 19660 4402 19672
rect 4617 19669 4629 19672
rect 4663 19669 4675 19703
rect 5108 19700 5136 19740
rect 5276 19740 5580 19768
rect 5276 19700 5304 19740
rect 5108 19672 5304 19700
rect 5552 19700 5580 19740
rect 5626 19728 5632 19780
rect 5684 19768 5690 19780
rect 5905 19771 5963 19777
rect 5905 19768 5917 19771
rect 5684 19740 5917 19768
rect 5684 19728 5690 19740
rect 5905 19737 5917 19740
rect 5951 19737 5963 19771
rect 5905 19731 5963 19737
rect 5810 19700 5816 19712
rect 5552 19672 5816 19700
rect 4617 19663 4675 19669
rect 5810 19660 5816 19672
rect 5868 19660 5874 19712
rect 5994 19660 6000 19712
rect 6052 19700 6058 19712
rect 6104 19700 6132 19808
rect 6641 19805 6653 19839
rect 6687 19836 6699 19839
rect 12526 19836 12532 19848
rect 6687 19808 12532 19836
rect 6687 19805 6699 19808
rect 6641 19799 6699 19805
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 6052 19672 6132 19700
rect 6457 19703 6515 19709
rect 6052 19660 6058 19672
rect 6457 19669 6469 19703
rect 6503 19700 6515 19703
rect 13998 19700 14004 19712
rect 6503 19672 14004 19700
rect 6503 19669 6515 19672
rect 6457 19663 6515 19669
rect 13998 19660 14004 19672
rect 14056 19660 14062 19712
rect 1104 19610 16836 19632
rect 1104 19558 4898 19610
rect 4950 19558 4962 19610
rect 5014 19558 5026 19610
rect 5078 19558 5090 19610
rect 5142 19558 5154 19610
rect 5206 19558 8846 19610
rect 8898 19558 8910 19610
rect 8962 19558 8974 19610
rect 9026 19558 9038 19610
rect 9090 19558 9102 19610
rect 9154 19558 12794 19610
rect 12846 19558 12858 19610
rect 12910 19558 12922 19610
rect 12974 19558 12986 19610
rect 13038 19558 13050 19610
rect 13102 19558 16836 19610
rect 1104 19536 16836 19558
rect 1397 19499 1455 19505
rect 1397 19465 1409 19499
rect 1443 19496 1455 19499
rect 1486 19496 1492 19508
rect 1443 19468 1492 19496
rect 1443 19465 1455 19468
rect 1397 19459 1455 19465
rect 1486 19456 1492 19468
rect 1544 19456 1550 19508
rect 3142 19496 3148 19508
rect 1596 19468 3148 19496
rect 1596 19428 1624 19468
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 3713 19499 3771 19505
rect 3713 19496 3725 19499
rect 3252 19468 3725 19496
rect 2590 19428 2596 19440
rect 1504 19400 1624 19428
rect 1872 19400 2596 19428
rect 1504 19372 1532 19400
rect 1486 19320 1492 19372
rect 1544 19320 1550 19372
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19329 1639 19363
rect 1581 19323 1639 19329
rect 1596 19292 1624 19323
rect 1670 19320 1676 19372
rect 1728 19360 1734 19372
rect 1728 19332 1773 19360
rect 1728 19320 1734 19332
rect 1872 19292 1900 19400
rect 2590 19388 2596 19400
rect 2648 19388 2654 19440
rect 2682 19388 2688 19440
rect 2740 19428 2746 19440
rect 3252 19428 3280 19468
rect 3713 19465 3725 19468
rect 3759 19465 3771 19499
rect 3713 19459 3771 19465
rect 4154 19456 4160 19508
rect 4212 19496 4218 19508
rect 4522 19496 4528 19508
rect 4212 19468 4528 19496
rect 4212 19456 4218 19468
rect 4522 19456 4528 19468
rect 4580 19456 4586 19508
rect 4908 19468 5396 19496
rect 3510 19428 3516 19440
rect 2740 19400 3280 19428
rect 3471 19400 3516 19428
rect 2740 19388 2746 19400
rect 3510 19388 3516 19400
rect 3568 19388 3574 19440
rect 4908 19437 4936 19468
rect 4893 19431 4951 19437
rect 4893 19397 4905 19431
rect 4939 19397 4951 19431
rect 4893 19391 4951 19397
rect 5123 19397 5181 19403
rect 1949 19363 2007 19369
rect 1949 19329 1961 19363
rect 1995 19360 2007 19363
rect 2314 19360 2320 19372
rect 1995 19332 2320 19360
rect 1995 19329 2007 19332
rect 1949 19323 2007 19329
rect 2314 19320 2320 19332
rect 2372 19320 2378 19372
rect 2774 19320 2780 19372
rect 2832 19360 2838 19372
rect 2961 19363 3019 19369
rect 2832 19332 2877 19360
rect 2832 19320 2838 19332
rect 2961 19329 2973 19363
rect 3007 19329 3019 19363
rect 5123 19363 5135 19397
rect 5169 19394 5181 19397
rect 5258 19394 5264 19440
rect 5169 19388 5264 19394
rect 5316 19388 5322 19440
rect 5169 19366 5304 19388
rect 5169 19363 5181 19366
rect 5123 19357 5181 19363
rect 5368 19360 5396 19468
rect 5534 19456 5540 19508
rect 5592 19496 5598 19508
rect 7101 19499 7159 19505
rect 7101 19496 7113 19499
rect 5592 19468 7113 19496
rect 5592 19456 5598 19468
rect 7101 19465 7113 19468
rect 7147 19465 7159 19499
rect 7101 19459 7159 19465
rect 6086 19388 6092 19440
rect 6144 19428 6150 19440
rect 6457 19431 6515 19437
rect 6457 19428 6469 19431
rect 6144 19400 6469 19428
rect 6144 19388 6150 19400
rect 6457 19397 6469 19400
rect 6503 19397 6515 19431
rect 15470 19428 15476 19440
rect 6457 19391 6515 19397
rect 6564 19400 15476 19428
rect 6564 19369 6592 19400
rect 15470 19388 15476 19400
rect 15528 19388 15534 19440
rect 6365 19363 6423 19369
rect 5368 19332 6316 19360
rect 2961 19323 3019 19329
rect 2038 19292 2044 19304
rect 1596 19264 1900 19292
rect 1999 19264 2044 19292
rect 2038 19252 2044 19264
rect 2096 19252 2102 19304
rect 2590 19252 2596 19304
rect 2648 19292 2654 19304
rect 2976 19292 3004 19323
rect 2648 19264 3004 19292
rect 3053 19295 3111 19301
rect 2648 19252 2654 19264
rect 3053 19261 3065 19295
rect 3099 19292 3111 19295
rect 5258 19292 5264 19304
rect 3099 19264 5264 19292
rect 3099 19261 3111 19264
rect 3053 19255 3111 19261
rect 5258 19252 5264 19264
rect 5316 19252 5322 19304
rect 3142 19184 3148 19236
rect 3200 19224 3206 19236
rect 3881 19227 3939 19233
rect 3881 19224 3893 19227
rect 3200 19196 3893 19224
rect 3200 19184 3206 19196
rect 3881 19193 3893 19196
rect 3927 19193 3939 19227
rect 5902 19224 5908 19236
rect 3881 19187 3939 19193
rect 5092 19196 5908 19224
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19156 3755 19159
rect 4798 19156 4804 19168
rect 3743 19128 4804 19156
rect 3743 19125 3755 19128
rect 3697 19119 3755 19125
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 5092 19165 5120 19196
rect 5902 19184 5908 19196
rect 5960 19184 5966 19236
rect 6288 19224 6316 19332
rect 6365 19329 6377 19363
rect 6411 19360 6423 19363
rect 6549 19363 6607 19369
rect 6411 19332 6500 19360
rect 6411 19329 6423 19332
rect 6365 19323 6423 19329
rect 6472 19292 6500 19332
rect 6549 19329 6561 19363
rect 6595 19329 6607 19363
rect 6549 19323 6607 19329
rect 6638 19320 6644 19372
rect 6696 19360 6702 19372
rect 7009 19363 7067 19369
rect 7009 19360 7021 19363
rect 6696 19332 7021 19360
rect 6696 19320 6702 19332
rect 7009 19329 7021 19332
rect 7055 19329 7067 19363
rect 10686 19360 10692 19372
rect 7009 19323 7067 19329
rect 7116 19332 10692 19360
rect 7116 19292 7144 19332
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 6472 19264 7144 19292
rect 7466 19224 7472 19236
rect 6288 19196 7472 19224
rect 7466 19184 7472 19196
rect 7524 19184 7530 19236
rect 17586 19224 17592 19236
rect 12406 19196 17592 19224
rect 5077 19159 5135 19165
rect 5077 19125 5089 19159
rect 5123 19125 5135 19159
rect 5077 19119 5135 19125
rect 5166 19116 5172 19168
rect 5224 19156 5230 19168
rect 5261 19159 5319 19165
rect 5261 19156 5273 19159
rect 5224 19128 5273 19156
rect 5224 19116 5230 19128
rect 5261 19125 5273 19128
rect 5307 19125 5319 19159
rect 5261 19119 5319 19125
rect 5810 19116 5816 19168
rect 5868 19156 5874 19168
rect 12406 19156 12434 19196
rect 17586 19184 17592 19196
rect 17644 19184 17650 19236
rect 5868 19128 12434 19156
rect 5868 19116 5874 19128
rect 1104 19066 16836 19088
rect 1104 19014 2924 19066
rect 2976 19014 2988 19066
rect 3040 19014 3052 19066
rect 3104 19014 3116 19066
rect 3168 19014 3180 19066
rect 3232 19014 6872 19066
rect 6924 19014 6936 19066
rect 6988 19014 7000 19066
rect 7052 19014 7064 19066
rect 7116 19014 7128 19066
rect 7180 19014 10820 19066
rect 10872 19014 10884 19066
rect 10936 19014 10948 19066
rect 11000 19014 11012 19066
rect 11064 19014 11076 19066
rect 11128 19014 14768 19066
rect 14820 19014 14832 19066
rect 14884 19014 14896 19066
rect 14948 19014 14960 19066
rect 15012 19014 15024 19066
rect 15076 19014 16836 19066
rect 1104 18992 16836 19014
rect 2501 18955 2559 18961
rect 2501 18921 2513 18955
rect 2547 18952 2559 18955
rect 2547 18924 3280 18952
rect 2547 18921 2559 18924
rect 2501 18915 2559 18921
rect 2774 18884 2780 18896
rect 2746 18844 2780 18884
rect 2832 18884 2838 18896
rect 3252 18884 3280 18924
rect 4706 18912 4712 18964
rect 4764 18952 4770 18964
rect 7193 18955 7251 18961
rect 4764 18924 6592 18952
rect 4764 18912 4770 18924
rect 3878 18884 3884 18896
rect 2832 18856 3188 18884
rect 3252 18856 3884 18884
rect 2832 18844 2838 18856
rect 2746 18816 2774 18844
rect 3050 18816 3056 18828
rect 1688 18788 2774 18816
rect 3011 18788 3056 18816
rect 1688 18757 1716 18788
rect 3050 18776 3056 18788
rect 3108 18776 3114 18828
rect 3160 18816 3188 18856
rect 3878 18844 3884 18856
rect 3936 18844 3942 18896
rect 3970 18844 3976 18896
rect 4028 18884 4034 18896
rect 4249 18887 4307 18893
rect 4249 18884 4261 18887
rect 4028 18856 4261 18884
rect 4028 18844 4034 18856
rect 4249 18853 4261 18856
rect 4295 18853 4307 18887
rect 6564 18884 6592 18924
rect 7193 18921 7205 18955
rect 7239 18952 7251 18955
rect 8294 18952 8300 18964
rect 7239 18924 8300 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 8294 18912 8300 18924
rect 8352 18912 8358 18964
rect 13906 18952 13912 18964
rect 8404 18924 13912 18952
rect 7745 18887 7803 18893
rect 7745 18884 7757 18887
rect 6564 18856 7757 18884
rect 4249 18847 4307 18853
rect 7745 18853 7757 18856
rect 7791 18853 7803 18887
rect 7745 18847 7803 18853
rect 3160 18788 5856 18816
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 1857 18751 1915 18757
rect 1857 18717 1869 18751
rect 1903 18717 1915 18751
rect 1857 18711 1915 18717
rect 1872 18612 1900 18711
rect 2314 18708 2320 18760
rect 2372 18748 2378 18760
rect 5445 18751 5503 18757
rect 5445 18748 5457 18751
rect 2372 18720 5457 18748
rect 2372 18708 2378 18720
rect 5445 18717 5457 18720
rect 5491 18717 5503 18751
rect 5718 18748 5724 18760
rect 5679 18720 5724 18748
rect 5445 18711 5503 18717
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 5828 18748 5856 18788
rect 6086 18776 6092 18828
rect 6144 18816 6150 18828
rect 8404 18816 8432 18924
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 8478 18844 8484 18896
rect 8536 18884 8542 18896
rect 13446 18884 13452 18896
rect 8536 18856 13452 18884
rect 8536 18844 8542 18856
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 6144 18788 8432 18816
rect 6144 18776 6150 18788
rect 6178 18748 6184 18760
rect 5828 18720 6184 18748
rect 6178 18708 6184 18720
rect 6236 18708 6242 18760
rect 6472 18757 6500 18788
rect 8754 18776 8760 18828
rect 8812 18816 8818 18828
rect 13814 18816 13820 18828
rect 8812 18788 13820 18816
rect 8812 18776 8818 18788
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18717 6515 18751
rect 6457 18711 6515 18717
rect 6546 18708 6552 18760
rect 6604 18748 6610 18760
rect 7098 18748 7104 18760
rect 6604 18720 6649 18748
rect 7059 18720 7104 18748
rect 6604 18708 6610 18720
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18748 7987 18751
rect 17034 18748 17040 18760
rect 7975 18720 17040 18748
rect 7975 18717 7987 18720
rect 7929 18711 7987 18717
rect 17034 18708 17040 18720
rect 17092 18708 17098 18760
rect 1949 18683 2007 18689
rect 1949 18649 1961 18683
rect 1995 18680 2007 18683
rect 2774 18680 2780 18692
rect 1995 18652 2780 18680
rect 1995 18649 2007 18652
rect 1949 18643 2007 18649
rect 2774 18640 2780 18652
rect 2832 18640 2838 18692
rect 3786 18680 3792 18692
rect 2884 18652 3792 18680
rect 2590 18612 2596 18624
rect 1872 18584 2596 18612
rect 2590 18572 2596 18584
rect 2648 18572 2654 18624
rect 2884 18621 2912 18652
rect 3786 18640 3792 18652
rect 3844 18640 3850 18692
rect 3973 18683 4031 18689
rect 3973 18649 3985 18683
rect 4019 18680 4031 18683
rect 4062 18680 4068 18692
rect 4019 18652 4068 18680
rect 4019 18649 4031 18652
rect 3973 18643 4031 18649
rect 4062 18640 4068 18652
rect 4120 18640 4126 18692
rect 5261 18683 5319 18689
rect 5261 18649 5273 18683
rect 5307 18680 5319 18683
rect 16850 18680 16856 18692
rect 5307 18652 16856 18680
rect 5307 18649 5319 18652
rect 5261 18643 5319 18649
rect 16850 18640 16856 18652
rect 16908 18640 16914 18692
rect 2869 18615 2927 18621
rect 2869 18581 2881 18615
rect 2915 18581 2927 18615
rect 2869 18575 2927 18581
rect 2961 18615 3019 18621
rect 2961 18581 2973 18615
rect 3007 18612 3019 18615
rect 3878 18612 3884 18624
rect 3007 18584 3884 18612
rect 3007 18581 3019 18584
rect 2961 18575 3019 18581
rect 3878 18572 3884 18584
rect 3936 18572 3942 18624
rect 4433 18615 4491 18621
rect 4433 18581 4445 18615
rect 4479 18612 4491 18615
rect 4522 18612 4528 18624
rect 4479 18584 4528 18612
rect 4479 18581 4491 18584
rect 4433 18575 4491 18581
rect 4522 18572 4528 18584
rect 4580 18572 4586 18624
rect 5629 18615 5687 18621
rect 5629 18581 5641 18615
rect 5675 18612 5687 18615
rect 5810 18612 5816 18624
rect 5675 18584 5816 18612
rect 5675 18581 5687 18584
rect 5629 18575 5687 18581
rect 5810 18572 5816 18584
rect 5868 18572 5874 18624
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 10778 18612 10784 18624
rect 8352 18584 10784 18612
rect 8352 18572 8358 18584
rect 10778 18572 10784 18584
rect 10836 18572 10842 18624
rect 1104 18522 16836 18544
rect 1104 18470 4898 18522
rect 4950 18470 4962 18522
rect 5014 18470 5026 18522
rect 5078 18470 5090 18522
rect 5142 18470 5154 18522
rect 5206 18470 8846 18522
rect 8898 18470 8910 18522
rect 8962 18470 8974 18522
rect 9026 18470 9038 18522
rect 9090 18470 9102 18522
rect 9154 18470 12794 18522
rect 12846 18470 12858 18522
rect 12910 18470 12922 18522
rect 12974 18470 12986 18522
rect 13038 18470 13050 18522
rect 13102 18470 16836 18522
rect 1104 18448 16836 18470
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 3234 18408 3240 18420
rect 2004 18380 3240 18408
rect 2004 18368 2010 18380
rect 3234 18368 3240 18380
rect 3292 18368 3298 18420
rect 3344 18380 4062 18408
rect 1302 18300 1308 18352
rect 1360 18340 1366 18352
rect 3344 18340 3372 18380
rect 1360 18312 3372 18340
rect 4034 18340 4062 18380
rect 6270 18368 6276 18420
rect 6328 18408 6334 18420
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 6328 18380 6561 18408
rect 6328 18368 6334 18380
rect 6549 18377 6561 18380
rect 6595 18377 6607 18411
rect 7466 18408 7472 18420
rect 7427 18380 7472 18408
rect 6549 18371 6607 18377
rect 7466 18368 7472 18380
rect 7524 18368 7530 18420
rect 8570 18368 8576 18420
rect 8628 18408 8634 18420
rect 8665 18411 8723 18417
rect 8665 18408 8677 18411
rect 8628 18380 8677 18408
rect 8628 18368 8634 18380
rect 8665 18377 8677 18380
rect 8711 18377 8723 18411
rect 8665 18371 8723 18377
rect 9030 18368 9036 18420
rect 9088 18408 9094 18420
rect 9306 18408 9312 18420
rect 9088 18380 9312 18408
rect 9088 18368 9094 18380
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 9490 18408 9496 18420
rect 9451 18380 9496 18408
rect 9490 18368 9496 18380
rect 9548 18368 9554 18420
rect 6365 18343 6423 18349
rect 4034 18312 5672 18340
rect 1360 18300 1366 18312
rect 1762 18232 1768 18284
rect 1820 18272 1826 18284
rect 2113 18275 2171 18281
rect 2113 18272 2125 18275
rect 1820 18244 2125 18272
rect 1820 18232 1826 18244
rect 2113 18241 2125 18244
rect 2159 18241 2171 18275
rect 2113 18235 2171 18241
rect 2866 18232 2872 18284
rect 2924 18272 2930 18284
rect 3694 18272 3700 18284
rect 2924 18244 3700 18272
rect 2924 18232 2930 18244
rect 3694 18232 3700 18244
rect 3752 18272 3758 18284
rect 5644 18281 5672 18312
rect 6365 18309 6377 18343
rect 6411 18340 6423 18343
rect 6454 18340 6460 18352
rect 6411 18312 6460 18340
rect 6411 18309 6423 18312
rect 6365 18303 6423 18309
rect 6454 18300 6460 18312
rect 6512 18300 6518 18352
rect 8113 18343 8171 18349
rect 8113 18309 8125 18343
rect 8159 18340 8171 18343
rect 9950 18340 9956 18352
rect 8159 18312 9956 18340
rect 8159 18309 8171 18312
rect 8113 18303 8171 18309
rect 9950 18300 9956 18312
rect 10008 18300 10014 18352
rect 4045 18275 4103 18281
rect 4045 18272 4057 18275
rect 3752 18244 4057 18272
rect 3752 18232 3758 18244
rect 4045 18241 4057 18244
rect 4091 18241 4103 18275
rect 4045 18235 4103 18241
rect 5629 18275 5687 18281
rect 5629 18241 5641 18275
rect 5675 18241 5687 18275
rect 5629 18235 5687 18241
rect 7190 18232 7196 18284
rect 7248 18272 7254 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 7248 18244 7389 18272
rect 7248 18232 7254 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 8018 18272 8024 18284
rect 7979 18244 8024 18272
rect 7377 18235 7435 18241
rect 8018 18232 8024 18244
rect 8076 18232 8082 18284
rect 8205 18275 8263 18281
rect 8205 18241 8217 18275
rect 8251 18272 8263 18275
rect 8294 18272 8300 18284
rect 8251 18244 8300 18272
rect 8251 18241 8263 18244
rect 8205 18235 8263 18241
rect 8294 18232 8300 18244
rect 8352 18232 8358 18284
rect 8849 18275 8907 18281
rect 8849 18241 8861 18275
rect 8895 18241 8907 18275
rect 8849 18235 8907 18241
rect 9309 18275 9367 18281
rect 9309 18241 9321 18275
rect 9355 18241 9367 18275
rect 9309 18235 9367 18241
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 16206 18272 16212 18284
rect 9539 18244 16212 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18173 1915 18207
rect 3786 18204 3792 18216
rect 3747 18176 3792 18204
rect 1857 18167 1915 18173
rect 1872 18068 1900 18167
rect 3786 18164 3792 18176
rect 3844 18164 3850 18216
rect 7466 18164 7472 18216
rect 7524 18204 7530 18216
rect 8864 18204 8892 18235
rect 7524 18176 8892 18204
rect 9324 18204 9352 18235
rect 16206 18232 16212 18244
rect 16264 18232 16270 18284
rect 11790 18204 11796 18216
rect 9324 18176 11796 18204
rect 7524 18164 7530 18176
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 3804 18136 3832 18164
rect 5813 18139 5871 18145
rect 5813 18136 5825 18139
rect 2792 18108 3832 18136
rect 4724 18108 5825 18136
rect 2792 18068 2820 18108
rect 1872 18040 2820 18068
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18068 3295 18071
rect 3418 18068 3424 18080
rect 3283 18040 3424 18068
rect 3283 18037 3295 18040
rect 3237 18031 3295 18037
rect 3418 18028 3424 18040
rect 3476 18028 3482 18080
rect 4062 18028 4068 18080
rect 4120 18068 4126 18080
rect 4724 18068 4752 18108
rect 5813 18105 5825 18108
rect 5859 18105 5871 18139
rect 5813 18099 5871 18105
rect 6733 18139 6791 18145
rect 6733 18105 6745 18139
rect 6779 18136 6791 18139
rect 12434 18136 12440 18148
rect 6779 18108 12440 18136
rect 6779 18105 6791 18108
rect 6733 18099 6791 18105
rect 12434 18096 12440 18108
rect 12492 18096 12498 18148
rect 5166 18068 5172 18080
rect 4120 18040 4752 18068
rect 5127 18040 5172 18068
rect 4120 18028 4126 18040
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6549 18071 6607 18077
rect 6549 18068 6561 18071
rect 6328 18040 6561 18068
rect 6328 18028 6334 18040
rect 6549 18037 6561 18040
rect 6595 18068 6607 18071
rect 8110 18068 8116 18080
rect 6595 18040 8116 18068
rect 6595 18037 6607 18040
rect 6549 18031 6607 18037
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 8754 18028 8760 18080
rect 8812 18068 8818 18080
rect 17126 18068 17132 18080
rect 8812 18040 17132 18068
rect 8812 18028 8818 18040
rect 17126 18028 17132 18040
rect 17184 18028 17190 18080
rect 1104 17978 16836 18000
rect 1104 17926 2924 17978
rect 2976 17926 2988 17978
rect 3040 17926 3052 17978
rect 3104 17926 3116 17978
rect 3168 17926 3180 17978
rect 3232 17926 6872 17978
rect 6924 17926 6936 17978
rect 6988 17926 7000 17978
rect 7052 17926 7064 17978
rect 7116 17926 7128 17978
rect 7180 17926 10820 17978
rect 10872 17926 10884 17978
rect 10936 17926 10948 17978
rect 11000 17926 11012 17978
rect 11064 17926 11076 17978
rect 11128 17926 14768 17978
rect 14820 17926 14832 17978
rect 14884 17926 14896 17978
rect 14948 17926 14960 17978
rect 15012 17926 15024 17978
rect 15076 17926 16836 17978
rect 1104 17904 16836 17926
rect 290 17824 296 17876
rect 348 17864 354 17876
rect 5629 17867 5687 17873
rect 5629 17864 5641 17867
rect 348 17836 5641 17864
rect 348 17824 354 17836
rect 5629 17833 5641 17836
rect 5675 17833 5687 17867
rect 5629 17827 5687 17833
rect 5718 17824 5724 17876
rect 5776 17864 5782 17876
rect 6270 17864 6276 17876
rect 5776 17836 6276 17864
rect 5776 17824 5782 17836
rect 6270 17824 6276 17836
rect 6328 17864 6334 17876
rect 6365 17867 6423 17873
rect 6365 17864 6377 17867
rect 6328 17836 6377 17864
rect 6328 17824 6334 17836
rect 6365 17833 6377 17836
rect 6411 17833 6423 17867
rect 6365 17827 6423 17833
rect 8941 17867 8999 17873
rect 8941 17833 8953 17867
rect 8987 17864 8999 17867
rect 9306 17864 9312 17876
rect 8987 17836 9312 17864
rect 8987 17833 8999 17836
rect 8941 17827 8999 17833
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 9416 17836 9628 17864
rect 3237 17799 3295 17805
rect 3237 17765 3249 17799
rect 3283 17765 3295 17799
rect 3237 17759 3295 17765
rect 3252 17728 3280 17759
rect 8018 17756 8024 17808
rect 8076 17796 8082 17808
rect 8205 17799 8263 17805
rect 8205 17796 8217 17799
rect 8076 17768 8217 17796
rect 8076 17756 8082 17768
rect 8205 17765 8217 17768
rect 8251 17765 8263 17799
rect 8205 17759 8263 17765
rect 8386 17756 8392 17808
rect 8444 17796 8450 17808
rect 9416 17796 9444 17836
rect 9600 17808 9628 17836
rect 10686 17824 10692 17876
rect 10744 17864 10750 17876
rect 15378 17864 15384 17876
rect 10744 17836 15384 17864
rect 10744 17824 10750 17836
rect 15378 17824 15384 17836
rect 15436 17824 15442 17876
rect 8444 17768 9444 17796
rect 8444 17756 8450 17768
rect 9582 17756 9588 17808
rect 9640 17756 9646 17808
rect 3252 17700 4384 17728
rect 1857 17663 1915 17669
rect 1857 17629 1869 17663
rect 1903 17660 1915 17663
rect 1946 17660 1952 17672
rect 1903 17632 1952 17660
rect 1903 17629 1915 17632
rect 1857 17623 1915 17629
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 4154 17660 4160 17672
rect 3528 17632 4160 17660
rect 1118 17552 1124 17604
rect 1176 17592 1182 17604
rect 2102 17595 2160 17601
rect 2102 17592 2114 17595
rect 1176 17564 2114 17592
rect 1176 17552 1182 17564
rect 2102 17561 2114 17564
rect 2148 17561 2160 17595
rect 2102 17555 2160 17561
rect 2117 17524 2145 17555
rect 2590 17552 2596 17604
rect 2648 17592 2654 17604
rect 3528 17592 3556 17632
rect 4154 17620 4160 17632
rect 4212 17660 4218 17672
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 4212 17632 4261 17660
rect 4212 17620 4218 17632
rect 4249 17629 4261 17632
rect 4295 17629 4307 17663
rect 4356 17660 4384 17700
rect 6086 17688 6092 17740
rect 6144 17728 6150 17740
rect 7466 17728 7472 17740
rect 6144 17700 7472 17728
rect 6144 17688 6150 17700
rect 7466 17688 7472 17700
rect 7524 17688 7530 17740
rect 8570 17688 8576 17740
rect 8628 17728 8634 17740
rect 9214 17728 9220 17740
rect 8628 17700 9220 17728
rect 8628 17688 8634 17700
rect 9214 17688 9220 17700
rect 9272 17688 9278 17740
rect 6641 17663 6699 17669
rect 4356 17632 4752 17660
rect 4249 17623 4307 17629
rect 4724 17604 4752 17632
rect 6641 17629 6653 17663
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17660 7343 17663
rect 7374 17660 7380 17672
rect 7331 17632 7380 17660
rect 7331 17629 7343 17632
rect 7285 17623 7343 17629
rect 2648 17564 3556 17592
rect 4494 17595 4552 17601
rect 2648 17552 2654 17564
rect 4494 17561 4506 17595
rect 4540 17561 4552 17595
rect 4494 17555 4552 17561
rect 3694 17524 3700 17536
rect 2117 17496 3700 17524
rect 3694 17484 3700 17496
rect 3752 17524 3758 17536
rect 4509 17524 4537 17555
rect 4706 17552 4712 17604
rect 4764 17552 4770 17604
rect 6181 17595 6239 17601
rect 6181 17561 6193 17595
rect 6227 17592 6239 17595
rect 6546 17592 6552 17604
rect 6227 17564 6552 17592
rect 6227 17561 6239 17564
rect 6181 17555 6239 17561
rect 6546 17552 6552 17564
rect 6604 17552 6610 17604
rect 3752 17496 4537 17524
rect 3752 17484 3758 17496
rect 5810 17484 5816 17536
rect 5868 17524 5874 17536
rect 6365 17527 6423 17533
rect 6365 17524 6377 17527
rect 5868 17496 6377 17524
rect 5868 17484 5874 17496
rect 6365 17493 6377 17496
rect 6411 17493 6423 17527
rect 6656 17524 6684 17623
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 7561 17663 7619 17669
rect 7561 17629 7573 17663
rect 7607 17660 7619 17663
rect 7742 17660 7748 17672
rect 7607 17632 7748 17660
rect 7607 17629 7619 17632
rect 7561 17623 7619 17629
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 8110 17620 8116 17672
rect 8168 17660 8174 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 8168 17632 8217 17660
rect 8168 17620 8174 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17629 8447 17663
rect 9122 17660 9128 17672
rect 8389 17623 8447 17629
rect 8588 17632 9128 17660
rect 7098 17592 7104 17604
rect 7059 17564 7104 17592
rect 7098 17552 7104 17564
rect 7156 17552 7162 17604
rect 7469 17595 7527 17601
rect 7469 17561 7481 17595
rect 7515 17592 7527 17595
rect 7834 17592 7840 17604
rect 7515 17564 7840 17592
rect 7515 17561 7527 17564
rect 7469 17555 7527 17561
rect 7834 17552 7840 17564
rect 7892 17552 7898 17604
rect 8404 17592 8432 17623
rect 8588 17604 8616 17632
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 9582 17620 9588 17672
rect 9640 17660 9646 17672
rect 9777 17663 9835 17669
rect 9640 17632 9685 17660
rect 9640 17620 9646 17632
rect 9777 17629 9789 17663
rect 9823 17660 9835 17663
rect 10134 17660 10140 17672
rect 9823 17632 10140 17660
rect 9823 17629 9835 17632
rect 9777 17623 9835 17629
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 8478 17592 8484 17604
rect 8404 17564 8484 17592
rect 8478 17552 8484 17564
rect 8536 17552 8542 17604
rect 8570 17552 8576 17604
rect 8628 17552 8634 17604
rect 9030 17552 9036 17604
rect 9088 17592 9094 17604
rect 9306 17592 9312 17604
rect 9088 17564 9312 17592
rect 9088 17552 9094 17564
rect 9306 17552 9312 17564
rect 9364 17552 9370 17604
rect 9490 17552 9496 17604
rect 9548 17592 9554 17604
rect 15654 17592 15660 17604
rect 9548 17564 15660 17592
rect 9548 17552 9554 17564
rect 15654 17552 15660 17564
rect 15712 17552 15718 17604
rect 8846 17524 8852 17536
rect 6656 17496 8852 17524
rect 6365 17487 6423 17493
rect 8846 17484 8852 17496
rect 8904 17484 8910 17536
rect 9769 17527 9827 17533
rect 9769 17493 9781 17527
rect 9815 17524 9827 17527
rect 10042 17524 10048 17536
rect 9815 17496 10048 17524
rect 9815 17493 9827 17496
rect 9769 17487 9827 17493
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 10226 17484 10232 17536
rect 10284 17524 10290 17536
rect 14458 17524 14464 17536
rect 10284 17496 14464 17524
rect 10284 17484 10290 17496
rect 14458 17484 14464 17496
rect 14516 17484 14522 17536
rect 1104 17434 16836 17456
rect 1104 17382 4898 17434
rect 4950 17382 4962 17434
rect 5014 17382 5026 17434
rect 5078 17382 5090 17434
rect 5142 17382 5154 17434
rect 5206 17382 8846 17434
rect 8898 17382 8910 17434
rect 8962 17382 8974 17434
rect 9026 17382 9038 17434
rect 9090 17382 9102 17434
rect 9154 17382 12794 17434
rect 12846 17382 12858 17434
rect 12910 17382 12922 17434
rect 12974 17382 12986 17434
rect 13038 17382 13050 17434
rect 13102 17382 16836 17434
rect 1104 17360 16836 17382
rect 3329 17323 3387 17329
rect 3329 17289 3341 17323
rect 3375 17320 3387 17323
rect 6454 17320 6460 17332
rect 3375 17292 6460 17320
rect 3375 17289 3387 17292
rect 3329 17283 3387 17289
rect 6454 17280 6460 17292
rect 6512 17280 6518 17332
rect 10226 17320 10232 17332
rect 6564 17292 10232 17320
rect 2130 17212 2136 17264
rect 2188 17252 2194 17264
rect 4034 17255 4092 17261
rect 4034 17252 4046 17255
rect 2188 17224 4046 17252
rect 2188 17212 2194 17224
rect 4034 17221 4046 17224
rect 4080 17221 4092 17255
rect 4034 17215 4092 17221
rect 1946 17184 1952 17196
rect 1907 17156 1952 17184
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 2216 17187 2274 17193
rect 2216 17153 2228 17187
rect 2262 17184 2274 17187
rect 2958 17184 2964 17196
rect 2262 17156 2964 17184
rect 2262 17153 2274 17156
rect 2216 17147 2274 17153
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 3786 17184 3792 17196
rect 3747 17156 3792 17184
rect 3786 17144 3792 17156
rect 3844 17144 3850 17196
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 5994 17184 6000 17196
rect 5859 17156 6000 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 5994 17144 6000 17156
rect 6052 17184 6058 17196
rect 6270 17184 6276 17196
rect 6052 17156 6276 17184
rect 6052 17144 6058 17156
rect 6270 17144 6276 17156
rect 6328 17144 6334 17196
rect 6564 17193 6592 17292
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 10686 17280 10692 17332
rect 10744 17320 10750 17332
rect 13630 17320 13636 17332
rect 10744 17292 13636 17320
rect 10744 17280 10750 17292
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 7650 17252 7656 17264
rect 6656 17224 7656 17252
rect 6656 17193 6684 17224
rect 7650 17212 7656 17224
rect 7708 17212 7714 17264
rect 7745 17255 7803 17261
rect 7745 17221 7757 17255
rect 7791 17252 7803 17255
rect 15746 17252 15752 17264
rect 7791 17224 15752 17252
rect 7791 17221 7803 17224
rect 7745 17215 7803 17221
rect 15746 17212 15752 17224
rect 15804 17212 15810 17264
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6641 17187 6699 17193
rect 6641 17153 6653 17187
rect 6687 17153 6699 17187
rect 6641 17147 6699 17153
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17184 7619 17187
rect 7834 17184 7840 17196
rect 7607 17156 7696 17184
rect 7795 17156 7840 17184
rect 7607 17153 7619 17156
rect 7561 17147 7619 17153
rect 6454 17076 6460 17128
rect 6512 17116 6518 17128
rect 6840 17116 6868 17147
rect 7374 17116 7380 17128
rect 6512 17088 6868 17116
rect 7335 17088 7380 17116
rect 6512 17076 6518 17088
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 5629 17051 5687 17057
rect 5629 17017 5641 17051
rect 5675 17048 5687 17051
rect 5718 17048 5724 17060
rect 5675 17020 5724 17048
rect 5675 17017 5687 17020
rect 5629 17011 5687 17017
rect 5718 17008 5724 17020
rect 5776 17008 5782 17060
rect 6733 17051 6791 17057
rect 6733 17017 6745 17051
rect 6779 17048 6791 17051
rect 7558 17048 7564 17060
rect 6779 17020 7564 17048
rect 6779 17017 6791 17020
rect 6733 17011 6791 17017
rect 7558 17008 7564 17020
rect 7616 17008 7622 17060
rect 7668 17048 7696 17156
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 7926 17144 7932 17196
rect 7984 17184 7990 17196
rect 8389 17187 8447 17193
rect 8389 17184 8401 17187
rect 7984 17156 8401 17184
rect 7984 17144 7990 17156
rect 8389 17153 8401 17156
rect 8435 17153 8447 17187
rect 9030 17184 9036 17196
rect 8943 17156 9036 17184
rect 8389 17147 8447 17153
rect 9030 17144 9036 17156
rect 9088 17184 9094 17196
rect 9674 17184 9680 17196
rect 9088 17156 9352 17184
rect 9635 17156 9680 17184
rect 9088 17144 9094 17156
rect 7742 17076 7748 17128
rect 7800 17116 7806 17128
rect 8570 17116 8576 17128
rect 7800 17088 8576 17116
rect 7800 17076 7806 17088
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 9324 17116 9352 17156
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 9858 17184 9864 17196
rect 9819 17156 9864 17184
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 10505 17187 10563 17193
rect 10505 17184 10517 17187
rect 10152 17156 10517 17184
rect 9876 17116 9904 17144
rect 9324 17088 9904 17116
rect 8018 17048 8024 17060
rect 7668 17020 8024 17048
rect 8018 17008 8024 17020
rect 8076 17008 8082 17060
rect 9398 17008 9404 17060
rect 9456 17048 9462 17060
rect 10152 17057 10180 17156
rect 10505 17153 10517 17156
rect 10551 17153 10563 17187
rect 10505 17147 10563 17153
rect 10318 17076 10324 17128
rect 10376 17116 10382 17128
rect 15102 17116 15108 17128
rect 10376 17088 15108 17116
rect 10376 17076 10382 17088
rect 15102 17076 15108 17088
rect 15160 17076 15166 17128
rect 10137 17051 10195 17057
rect 10137 17048 10149 17051
rect 9456 17020 10149 17048
rect 9456 17008 9462 17020
rect 10137 17017 10149 17020
rect 10183 17017 10195 17051
rect 10137 17011 10195 17017
rect 10689 17051 10747 17057
rect 10689 17017 10701 17051
rect 10735 17048 10747 17051
rect 16758 17048 16764 17060
rect 10735 17020 16764 17048
rect 10735 17017 10747 17020
rect 10689 17011 10747 17017
rect 16758 17008 16764 17020
rect 16816 17008 16822 17060
rect 4430 16940 4436 16992
rect 4488 16980 4494 16992
rect 5169 16983 5227 16989
rect 5169 16980 5181 16983
rect 4488 16952 5181 16980
rect 4488 16940 4494 16952
rect 5169 16949 5181 16952
rect 5215 16949 5227 16983
rect 5169 16943 5227 16949
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 6365 16983 6423 16989
rect 6365 16980 6377 16983
rect 6052 16952 6377 16980
rect 6052 16940 6058 16952
rect 6365 16949 6377 16952
rect 6411 16949 6423 16983
rect 6365 16943 6423 16949
rect 6638 16940 6644 16992
rect 6696 16980 6702 16992
rect 8481 16983 8539 16989
rect 8481 16980 8493 16983
rect 6696 16952 8493 16980
rect 6696 16940 6702 16952
rect 8481 16949 8493 16952
rect 8527 16949 8539 16983
rect 8481 16943 8539 16949
rect 9125 16983 9183 16989
rect 9125 16949 9137 16983
rect 9171 16980 9183 16983
rect 9674 16980 9680 16992
rect 9171 16952 9680 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 9769 16983 9827 16989
rect 9769 16949 9781 16983
rect 9815 16980 9827 16983
rect 10502 16980 10508 16992
rect 9815 16952 10508 16980
rect 9815 16949 9827 16952
rect 9769 16943 9827 16949
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 10594 16940 10600 16992
rect 10652 16980 10658 16992
rect 14274 16980 14280 16992
rect 10652 16952 14280 16980
rect 10652 16940 10658 16952
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 1104 16890 16836 16912
rect 1104 16838 2924 16890
rect 2976 16838 2988 16890
rect 3040 16838 3052 16890
rect 3104 16838 3116 16890
rect 3168 16838 3180 16890
rect 3232 16838 6872 16890
rect 6924 16838 6936 16890
rect 6988 16838 7000 16890
rect 7052 16838 7064 16890
rect 7116 16838 7128 16890
rect 7180 16838 10820 16890
rect 10872 16838 10884 16890
rect 10936 16838 10948 16890
rect 11000 16838 11012 16890
rect 11064 16838 11076 16890
rect 11128 16838 14768 16890
rect 14820 16838 14832 16890
rect 14884 16838 14896 16890
rect 14948 16838 14960 16890
rect 15012 16838 15024 16890
rect 15076 16838 16836 16890
rect 1104 16816 16836 16838
rect 842 16736 848 16788
rect 900 16776 906 16788
rect 900 16748 2903 16776
rect 900 16736 906 16748
rect 2875 16640 2903 16748
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 6549 16779 6607 16785
rect 6549 16776 6561 16779
rect 6236 16748 6561 16776
rect 6236 16736 6242 16748
rect 6549 16745 6561 16748
rect 6595 16745 6607 16779
rect 6549 16739 6607 16745
rect 7742 16736 7748 16788
rect 7800 16776 7806 16788
rect 8018 16776 8024 16788
rect 7800 16748 8024 16776
rect 7800 16736 7806 16748
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 9490 16776 9496 16788
rect 8352 16748 9496 16776
rect 8352 16736 8358 16748
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 10318 16776 10324 16788
rect 9824 16748 10324 16776
rect 9824 16736 9830 16748
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 10597 16779 10655 16785
rect 10597 16745 10609 16779
rect 10643 16745 10655 16779
rect 10597 16739 10655 16745
rect 5442 16668 5448 16720
rect 5500 16708 5506 16720
rect 5500 16680 8800 16708
rect 5500 16668 5506 16680
rect 2875 16612 6316 16640
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16572 1915 16575
rect 2590 16572 2596 16584
rect 1903 16544 2596 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 2590 16532 2596 16544
rect 2648 16532 2654 16584
rect 4522 16532 4528 16584
rect 4580 16572 4586 16584
rect 6288 16572 6316 16612
rect 6362 16600 6368 16652
rect 6420 16640 6426 16652
rect 8772 16640 8800 16680
rect 8938 16668 8944 16720
rect 8996 16708 9002 16720
rect 10612 16708 10640 16739
rect 10778 16736 10784 16788
rect 10836 16776 10842 16788
rect 16574 16776 16580 16788
rect 10836 16748 16580 16776
rect 10836 16736 10842 16748
rect 16574 16736 16580 16748
rect 16632 16736 16638 16788
rect 8996 16680 10640 16708
rect 11517 16711 11575 16717
rect 8996 16668 9002 16680
rect 11517 16677 11529 16711
rect 11563 16677 11575 16711
rect 11517 16671 11575 16677
rect 10594 16640 10600 16652
rect 6420 16612 8708 16640
rect 8772 16612 10600 16640
rect 6420 16600 6426 16612
rect 7929 16575 7987 16581
rect 7929 16572 7941 16575
rect 4580 16544 4625 16572
rect 6288 16544 7941 16572
rect 4580 16532 4586 16544
rect 7929 16541 7941 16544
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16572 8171 16575
rect 8294 16572 8300 16584
rect 8159 16544 8300 16572
rect 8159 16541 8171 16544
rect 8113 16535 8171 16541
rect 8294 16532 8300 16544
rect 8352 16532 8358 16584
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16572 8447 16575
rect 8570 16572 8576 16584
rect 8435 16544 8576 16572
rect 8435 16541 8447 16544
rect 8389 16535 8447 16541
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 8680 16582 8708 16612
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 8680 16572 8800 16582
rect 8938 16572 8944 16584
rect 8680 16554 8944 16572
rect 8772 16544 8944 16554
rect 8938 16532 8944 16544
rect 8996 16532 9002 16584
rect 9122 16532 9128 16584
rect 9180 16572 9186 16584
rect 11532 16572 11560 16671
rect 11698 16572 11704 16584
rect 9180 16544 11560 16572
rect 11659 16544 11704 16572
rect 9180 16532 9186 16544
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 1762 16464 1768 16516
rect 1820 16504 1826 16516
rect 2102 16507 2160 16513
rect 2102 16504 2114 16507
rect 1820 16476 2114 16504
rect 1820 16464 1826 16476
rect 2102 16473 2114 16476
rect 2148 16473 2160 16507
rect 2102 16467 2160 16473
rect 2424 16476 3464 16504
rect 750 16396 756 16448
rect 808 16436 814 16448
rect 1486 16436 1492 16448
rect 808 16408 1492 16436
rect 808 16396 814 16408
rect 1486 16396 1492 16408
rect 1544 16436 1550 16448
rect 2424 16436 2452 16476
rect 1544 16408 2452 16436
rect 3237 16439 3295 16445
rect 1544 16396 1550 16408
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 3326 16436 3332 16448
rect 3283 16408 3332 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 3326 16396 3332 16408
rect 3384 16396 3390 16448
rect 3436 16436 3464 16476
rect 4062 16464 4068 16516
rect 4120 16504 4126 16516
rect 4249 16507 4307 16513
rect 4249 16504 4261 16507
rect 4120 16476 4261 16504
rect 4120 16464 4126 16476
rect 4249 16473 4261 16476
rect 4295 16473 4307 16507
rect 4249 16467 4307 16473
rect 5261 16507 5319 16513
rect 5261 16473 5273 16507
rect 5307 16504 5319 16507
rect 7098 16504 7104 16516
rect 5307 16476 7104 16504
rect 5307 16473 5319 16476
rect 5261 16467 5319 16473
rect 7098 16464 7104 16476
rect 7156 16464 7162 16516
rect 4433 16439 4491 16445
rect 4433 16436 4445 16439
rect 3436 16408 4445 16436
rect 4433 16405 4445 16408
rect 4479 16405 4491 16439
rect 4614 16436 4620 16448
rect 4575 16408 4620 16436
rect 4433 16399 4491 16405
rect 4614 16396 4620 16408
rect 4672 16396 4678 16448
rect 4798 16436 4804 16448
rect 4759 16408 4804 16436
rect 4798 16396 4804 16408
rect 4856 16396 4862 16448
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 6362 16436 6368 16448
rect 5592 16408 6368 16436
rect 5592 16396 5598 16408
rect 6362 16396 6368 16408
rect 6420 16396 6426 16448
rect 6822 16396 6828 16448
rect 6880 16436 6886 16448
rect 7282 16436 7288 16448
rect 6880 16408 7288 16436
rect 6880 16396 6886 16408
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 7374 16396 7380 16448
rect 7432 16436 7438 16448
rect 8202 16436 8208 16448
rect 7432 16408 8208 16436
rect 7432 16396 7438 16408
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 8297 16439 8355 16445
rect 8297 16405 8309 16439
rect 8343 16436 8355 16439
rect 8478 16436 8484 16448
rect 8343 16408 8484 16436
rect 8343 16405 8355 16408
rect 8297 16399 8355 16405
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 8588 16436 8616 16532
rect 8662 16464 8668 16516
rect 8720 16504 8726 16516
rect 9214 16504 9220 16516
rect 8720 16476 9220 16504
rect 8720 16464 8726 16476
rect 9214 16464 9220 16476
rect 9272 16464 9278 16516
rect 9309 16507 9367 16513
rect 9309 16473 9321 16507
rect 9355 16504 9367 16507
rect 14550 16504 14556 16516
rect 9355 16476 11376 16504
rect 9355 16473 9367 16476
rect 9309 16467 9367 16473
rect 9674 16436 9680 16448
rect 8588 16408 9680 16436
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 9858 16396 9864 16448
rect 9916 16436 9922 16448
rect 10870 16436 10876 16448
rect 9916 16408 10876 16436
rect 9916 16396 9922 16408
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11348 16436 11376 16476
rect 12406 16476 14556 16504
rect 12406 16436 12434 16476
rect 14550 16464 14556 16476
rect 14608 16464 14614 16516
rect 11348 16408 12434 16436
rect 1104 16346 16836 16368
rect 1104 16294 4898 16346
rect 4950 16294 4962 16346
rect 5014 16294 5026 16346
rect 5078 16294 5090 16346
rect 5142 16294 5154 16346
rect 5206 16294 8846 16346
rect 8898 16294 8910 16346
rect 8962 16294 8974 16346
rect 9026 16294 9038 16346
rect 9090 16294 9102 16346
rect 9154 16294 12794 16346
rect 12846 16294 12858 16346
rect 12910 16294 12922 16346
rect 12974 16294 12986 16346
rect 13038 16294 13050 16346
rect 13102 16294 16836 16346
rect 1104 16272 16836 16294
rect 1397 16235 1455 16241
rect 1397 16201 1409 16235
rect 1443 16232 1455 16235
rect 2222 16232 2228 16244
rect 1443 16204 2228 16232
rect 1443 16201 1455 16204
rect 1397 16195 1455 16201
rect 2222 16192 2228 16204
rect 2280 16192 2286 16244
rect 2406 16192 2412 16244
rect 2464 16232 2470 16244
rect 2682 16232 2688 16244
rect 2464 16204 2688 16232
rect 2464 16192 2470 16204
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 8018 16232 8024 16244
rect 4715 16204 8024 16232
rect 2498 16164 2504 16176
rect 1688 16136 2504 16164
rect 1210 16056 1216 16108
rect 1268 16096 1274 16108
rect 1688 16105 1716 16136
rect 2498 16124 2504 16136
rect 2556 16124 2562 16176
rect 2866 16173 2872 16176
rect 2860 16164 2872 16173
rect 2827 16136 2872 16164
rect 2860 16127 2872 16136
rect 2866 16124 2872 16127
rect 2924 16124 2930 16176
rect 3970 16124 3976 16176
rect 4028 16164 4034 16176
rect 4522 16164 4528 16176
rect 4028 16136 4528 16164
rect 4028 16124 4034 16136
rect 4522 16124 4528 16136
rect 4580 16124 4586 16176
rect 4715 16173 4743 16204
rect 8018 16192 8024 16204
rect 8076 16192 8082 16244
rect 8294 16232 8300 16244
rect 8128 16204 8300 16232
rect 4700 16167 4758 16173
rect 4700 16133 4712 16167
rect 4746 16133 4758 16167
rect 4700 16127 4758 16133
rect 5902 16124 5908 16176
rect 5960 16164 5966 16176
rect 6917 16167 6975 16173
rect 5960 16136 6224 16164
rect 5960 16124 5966 16136
rect 6196 16108 6224 16136
rect 6917 16133 6929 16167
rect 6963 16164 6975 16167
rect 8128 16164 8156 16204
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 8754 16232 8760 16244
rect 8404 16204 8760 16232
rect 6963 16136 8156 16164
rect 8201 16167 8259 16173
rect 6963 16133 6975 16136
rect 6917 16127 6975 16133
rect 8201 16133 8213 16167
rect 8247 16164 8259 16167
rect 8404 16164 8432 16204
rect 8754 16192 8760 16204
rect 8812 16192 8818 16244
rect 9766 16232 9772 16244
rect 8864 16204 9772 16232
rect 8247 16136 8432 16164
rect 8247 16133 8259 16136
rect 8201 16127 8259 16133
rect 8478 16124 8484 16176
rect 8536 16164 8542 16176
rect 8864 16164 8892 16204
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 10594 16192 10600 16244
rect 10652 16232 10658 16244
rect 10652 16204 12112 16232
rect 10652 16192 10658 16204
rect 8536 16136 8892 16164
rect 8536 16124 8542 16136
rect 9398 16124 9404 16176
rect 9456 16164 9462 16176
rect 9456 16136 9996 16164
rect 9456 16124 9462 16136
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1268 16068 1685 16096
rect 1268 16056 1274 16068
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 2222 16096 2228 16108
rect 1811 16068 2228 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 6178 16056 6184 16108
rect 6236 16096 6242 16108
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 6236 16068 6377 16096
rect 6236 16056 6242 16068
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6638 16096 6644 16108
rect 6599 16068 6644 16096
rect 6365 16059 6423 16065
rect 6638 16056 6644 16068
rect 6696 16056 6702 16108
rect 6730 16056 6736 16108
rect 6788 16096 6794 16108
rect 7190 16096 7196 16108
rect 6788 16068 7196 16096
rect 6788 16056 6794 16068
rect 7190 16056 7196 16068
rect 7248 16056 7254 16108
rect 7926 16096 7932 16108
rect 7887 16068 7932 16096
rect 7926 16056 7932 16068
rect 7984 16056 7990 16108
rect 8110 16096 8116 16108
rect 8071 16068 8116 16096
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 8294 16096 8300 16108
rect 8255 16068 8300 16096
rect 8294 16056 8300 16068
rect 8352 16096 8358 16108
rect 9582 16096 9588 16108
rect 8352 16068 9588 16096
rect 8352 16056 8358 16068
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16065 9735 16099
rect 9858 16096 9864 16108
rect 9819 16068 9864 16096
rect 9677 16059 9735 16065
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 1854 16028 1860 16040
rect 1815 16000 1860 16028
rect 1854 15988 1860 16000
rect 1912 15988 1918 16040
rect 2590 16028 2596 16040
rect 2551 16000 2596 16028
rect 2590 15988 2596 16000
rect 2648 15988 2654 16040
rect 4433 16031 4491 16037
rect 4433 15997 4445 16031
rect 4479 15997 4491 16031
rect 9306 16028 9312 16040
rect 4433 15991 4491 15997
rect 6564 16000 9312 16028
rect 3694 15852 3700 15904
rect 3752 15892 3758 15904
rect 3973 15895 4031 15901
rect 3973 15892 3985 15895
rect 3752 15864 3985 15892
rect 3752 15852 3758 15864
rect 3973 15861 3985 15864
rect 4019 15861 4031 15895
rect 4448 15892 4476 15991
rect 5902 15920 5908 15972
rect 5960 15960 5966 15972
rect 6564 15960 6592 16000
rect 9306 15988 9312 16000
rect 9364 15988 9370 16040
rect 9692 16028 9720 16059
rect 9858 16056 9864 16068
rect 9916 16056 9922 16108
rect 9968 16105 9996 16136
rect 10226 16124 10232 16176
rect 10284 16164 10290 16176
rect 10781 16167 10839 16173
rect 10781 16164 10793 16167
rect 10284 16136 10793 16164
rect 10284 16124 10290 16136
rect 10781 16133 10793 16136
rect 10827 16133 10839 16167
rect 12084 16164 12112 16204
rect 12158 16192 12164 16244
rect 12216 16232 12222 16244
rect 15289 16235 15347 16241
rect 15289 16232 15301 16235
rect 12216 16204 15301 16232
rect 12216 16192 12222 16204
rect 15289 16201 15301 16204
rect 15335 16201 15347 16235
rect 15289 16195 15347 16201
rect 14090 16164 14096 16176
rect 12084 16136 14096 16164
rect 10781 16127 10839 16133
rect 14090 16124 14096 16136
rect 14148 16124 14154 16176
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16065 10011 16099
rect 10594 16096 10600 16108
rect 10555 16068 10600 16096
rect 9953 16059 10011 16065
rect 10594 16056 10600 16068
rect 10652 16056 10658 16108
rect 10870 16096 10876 16108
rect 10783 16068 10876 16096
rect 10870 16056 10876 16068
rect 10928 16096 10934 16108
rect 11606 16096 11612 16108
rect 10928 16068 11612 16096
rect 10928 16056 10934 16068
rect 11606 16056 11612 16068
rect 11664 16056 11670 16108
rect 11701 16099 11759 16105
rect 11701 16065 11713 16099
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11238 16028 11244 16040
rect 9692 16000 11244 16028
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 11716 16028 11744 16059
rect 11882 16056 11888 16108
rect 11940 16096 11946 16108
rect 12345 16099 12403 16105
rect 12345 16096 12357 16099
rect 11940 16068 12357 16096
rect 11940 16056 11946 16068
rect 12345 16065 12357 16068
rect 12391 16065 12403 16099
rect 12345 16059 12403 16065
rect 15286 16056 15292 16108
rect 15344 16096 15350 16108
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15344 16068 15485 16096
rect 15344 16056 15350 16068
rect 15473 16065 15485 16068
rect 15519 16096 15531 16099
rect 16482 16096 16488 16108
rect 15519 16068 16488 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 11716 16000 15332 16028
rect 15304 15972 15332 16000
rect 5960 15932 6592 15960
rect 5960 15920 5966 15932
rect 7098 15920 7104 15972
rect 7156 15960 7162 15972
rect 8662 15960 8668 15972
rect 7156 15932 8668 15960
rect 7156 15920 7162 15932
rect 8662 15920 8668 15932
rect 8720 15920 8726 15972
rect 8846 15920 8852 15972
rect 8904 15960 8910 15972
rect 8904 15932 9820 15960
rect 8904 15920 8910 15932
rect 5718 15892 5724 15904
rect 4448 15864 5724 15892
rect 3973 15855 4031 15861
rect 5718 15852 5724 15864
rect 5776 15852 5782 15904
rect 5813 15895 5871 15901
rect 5813 15861 5825 15895
rect 5859 15892 5871 15895
rect 6362 15892 6368 15904
rect 5859 15864 6368 15892
rect 5859 15861 5871 15864
rect 5813 15855 5871 15861
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 6638 15852 6644 15904
rect 6696 15892 6702 15904
rect 6822 15892 6828 15904
rect 6696 15864 6828 15892
rect 6696 15852 6702 15864
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 6914 15852 6920 15904
rect 6972 15892 6978 15904
rect 8294 15892 8300 15904
rect 6972 15864 8300 15892
rect 6972 15852 6978 15864
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 8481 15895 8539 15901
rect 8481 15861 8493 15895
rect 8527 15892 8539 15895
rect 8754 15892 8760 15904
rect 8527 15864 8760 15892
rect 8527 15861 8539 15864
rect 8481 15855 8539 15861
rect 8754 15852 8760 15864
rect 8812 15852 8818 15904
rect 9493 15895 9551 15901
rect 9493 15861 9505 15895
rect 9539 15892 9551 15895
rect 9582 15892 9588 15904
rect 9539 15864 9588 15892
rect 9539 15861 9551 15864
rect 9493 15855 9551 15861
rect 9582 15852 9588 15864
rect 9640 15852 9646 15904
rect 9792 15892 9820 15932
rect 9858 15920 9864 15972
rect 9916 15960 9922 15972
rect 12618 15960 12624 15972
rect 9916 15932 12624 15960
rect 9916 15920 9922 15932
rect 12618 15920 12624 15932
rect 12676 15920 12682 15972
rect 15286 15920 15292 15972
rect 15344 15920 15350 15972
rect 9950 15892 9956 15904
rect 9792 15864 9956 15892
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10413 15895 10471 15901
rect 10413 15861 10425 15895
rect 10459 15892 10471 15895
rect 10686 15892 10692 15904
rect 10459 15864 10692 15892
rect 10459 15861 10471 15864
rect 10413 15855 10471 15861
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 10778 15852 10784 15904
rect 10836 15892 10842 15904
rect 11330 15892 11336 15904
rect 10836 15864 11336 15892
rect 10836 15852 10842 15864
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 11514 15892 11520 15904
rect 11475 15864 11520 15892
rect 11514 15852 11520 15864
rect 11572 15852 11578 15904
rect 11698 15852 11704 15904
rect 11756 15892 11762 15904
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 11756 15864 12173 15892
rect 11756 15852 11762 15864
rect 12161 15861 12173 15864
rect 12207 15861 12219 15895
rect 12161 15855 12219 15861
rect 1104 15802 16836 15824
rect 1104 15750 2924 15802
rect 2976 15750 2988 15802
rect 3040 15750 3052 15802
rect 3104 15750 3116 15802
rect 3168 15750 3180 15802
rect 3232 15750 6872 15802
rect 6924 15750 6936 15802
rect 6988 15750 7000 15802
rect 7052 15750 7064 15802
rect 7116 15750 7128 15802
rect 7180 15750 10820 15802
rect 10872 15750 10884 15802
rect 10936 15750 10948 15802
rect 11000 15750 11012 15802
rect 11064 15750 11076 15802
rect 11128 15750 14768 15802
rect 14820 15750 14832 15802
rect 14884 15750 14896 15802
rect 14948 15750 14960 15802
rect 15012 15750 15024 15802
rect 15076 15750 16836 15802
rect 1104 15728 16836 15750
rect 2130 15688 2136 15700
rect 1412 15660 2136 15688
rect 1412 15632 1440 15660
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 3970 15688 3976 15700
rect 3931 15660 3976 15688
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 4801 15691 4859 15697
rect 4801 15657 4813 15691
rect 4847 15688 4859 15691
rect 5626 15688 5632 15700
rect 4847 15660 5632 15688
rect 4847 15657 4859 15660
rect 4801 15651 4859 15657
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 6546 15688 6552 15700
rect 6507 15660 6552 15688
rect 6546 15648 6552 15660
rect 6604 15648 6610 15700
rect 12158 15688 12164 15700
rect 6886 15660 12164 15688
rect 1394 15580 1400 15632
rect 1452 15580 1458 15632
rect 2590 15620 2596 15632
rect 2424 15592 2596 15620
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15484 1455 15487
rect 2424 15484 2452 15592
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 3786 15580 3792 15632
rect 3844 15620 3850 15632
rect 4154 15620 4160 15632
rect 3844 15592 4160 15620
rect 3844 15580 3850 15592
rect 4154 15580 4160 15592
rect 4212 15580 4218 15632
rect 2498 15512 2504 15564
rect 2556 15552 2562 15564
rect 6886 15552 6914 15660
rect 12158 15648 12164 15660
rect 12216 15648 12222 15700
rect 13078 15688 13084 15700
rect 13039 15660 13084 15688
rect 13078 15648 13084 15660
rect 13136 15648 13142 15700
rect 14550 15688 14556 15700
rect 14511 15660 14556 15688
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 7742 15580 7748 15632
rect 7800 15620 7806 15632
rect 10962 15629 10968 15632
rect 10919 15623 10968 15629
rect 7800 15592 10272 15620
rect 7800 15580 7806 15592
rect 2556 15524 6914 15552
rect 8113 15555 8171 15561
rect 2556 15512 2562 15524
rect 8113 15521 8125 15555
rect 8159 15552 8171 15555
rect 8294 15552 8300 15564
rect 8159 15524 8300 15552
rect 8159 15521 8171 15524
rect 8113 15515 8171 15521
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 9490 15512 9496 15564
rect 9548 15552 9554 15564
rect 9548 15524 10088 15552
rect 9548 15512 9554 15524
rect 10060 15496 10088 15524
rect 1443 15456 2452 15484
rect 1443 15453 1455 15456
rect 1397 15447 1455 15453
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 3973 15487 4031 15493
rect 3973 15484 3985 15487
rect 3844 15456 3985 15484
rect 3844 15444 3850 15456
rect 3973 15453 3985 15456
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4617 15487 4675 15493
rect 4203 15456 4568 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 1642 15419 1700 15425
rect 1642 15416 1654 15419
rect 1412 15388 1654 15416
rect 1412 15360 1440 15388
rect 1642 15385 1654 15388
rect 1688 15385 1700 15419
rect 1642 15379 1700 15385
rect 2314 15376 2320 15428
rect 2372 15416 2378 15428
rect 4338 15416 4344 15428
rect 2372 15388 4344 15416
rect 2372 15376 2378 15388
rect 4338 15376 4344 15388
rect 4396 15376 4402 15428
rect 1394 15308 1400 15360
rect 1452 15308 1458 15360
rect 2777 15351 2835 15357
rect 2777 15317 2789 15351
rect 2823 15348 2835 15351
rect 3970 15348 3976 15360
rect 2823 15320 3976 15348
rect 2823 15317 2835 15320
rect 2777 15311 2835 15317
rect 3970 15308 3976 15320
rect 4028 15308 4034 15360
rect 4540 15348 4568 15456
rect 4617 15453 4629 15487
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15484 5319 15487
rect 5534 15484 5540 15496
rect 5307 15456 5540 15484
rect 5307 15453 5319 15456
rect 5261 15447 5319 15453
rect 4632 15416 4660 15447
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15484 7895 15487
rect 8478 15484 8484 15496
rect 7883 15456 8484 15484
rect 7883 15453 7895 15456
rect 7837 15447 7895 15453
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 9030 15444 9036 15496
rect 9088 15484 9094 15496
rect 9144 15487 9202 15493
rect 9144 15484 9156 15487
rect 9088 15456 9156 15484
rect 9088 15444 9094 15456
rect 9144 15453 9156 15456
rect 9190 15453 9202 15487
rect 9144 15447 9202 15453
rect 9398 15444 9404 15496
rect 9456 15484 9462 15496
rect 10042 15484 10048 15496
rect 9456 15456 9501 15484
rect 10003 15456 10048 15484
rect 9456 15444 9462 15456
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 10244 15493 10272 15592
rect 10919 15589 10931 15623
rect 10965 15589 10968 15623
rect 10919 15583 10968 15589
rect 10962 15580 10968 15583
rect 11020 15580 11026 15632
rect 11330 15580 11336 15632
rect 11388 15620 11394 15632
rect 12345 15623 12403 15629
rect 12345 15620 12357 15623
rect 11388 15592 12357 15620
rect 11388 15580 11394 15592
rect 12345 15589 12357 15592
rect 12391 15589 12403 15623
rect 12345 15583 12403 15589
rect 12526 15580 12532 15632
rect 12584 15620 12590 15632
rect 12584 15592 13124 15620
rect 12584 15580 12590 15592
rect 11054 15552 11060 15564
rect 11015 15524 11060 15552
rect 11054 15512 11060 15524
rect 11112 15512 11118 15564
rect 11149 15555 11207 15561
rect 11149 15521 11161 15555
rect 11195 15552 11207 15555
rect 12250 15552 12256 15564
rect 11195 15524 12256 15552
rect 11195 15521 11207 15524
rect 11149 15515 11207 15521
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 12894 15552 12900 15564
rect 12452 15524 12900 15552
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10318 15444 10324 15496
rect 10376 15484 10382 15496
rect 10778 15484 10784 15496
rect 10376 15456 10421 15484
rect 10739 15456 10784 15484
rect 10376 15444 10382 15456
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15484 11299 15487
rect 11422 15484 11428 15496
rect 11287 15456 11428 15484
rect 11287 15453 11299 15456
rect 11241 15447 11299 15453
rect 4632 15388 10456 15416
rect 10060 15360 10088 15388
rect 5074 15348 5080 15360
rect 4540 15320 5080 15348
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 6086 15308 6092 15360
rect 6144 15348 6150 15360
rect 7469 15351 7527 15357
rect 7469 15348 7481 15351
rect 6144 15320 7481 15348
rect 6144 15308 6150 15320
rect 7469 15317 7481 15320
rect 7515 15317 7527 15351
rect 7469 15311 7527 15317
rect 7929 15351 7987 15357
rect 7929 15317 7941 15351
rect 7975 15348 7987 15351
rect 8662 15348 8668 15360
rect 7975 15320 8668 15348
rect 7975 15317 7987 15320
rect 7929 15311 7987 15317
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 8938 15348 8944 15360
rect 8899 15320 8944 15348
rect 8938 15308 8944 15320
rect 8996 15308 9002 15360
rect 9214 15308 9220 15360
rect 9272 15348 9278 15360
rect 9309 15351 9367 15357
rect 9309 15348 9321 15351
rect 9272 15320 9321 15348
rect 9272 15308 9278 15320
rect 9309 15317 9321 15320
rect 9355 15317 9367 15351
rect 9858 15348 9864 15360
rect 9819 15320 9864 15348
rect 9309 15311 9367 15317
rect 9858 15308 9864 15320
rect 9916 15308 9922 15360
rect 10042 15308 10048 15360
rect 10100 15308 10106 15360
rect 10428 15348 10456 15388
rect 10594 15376 10600 15428
rect 10652 15416 10658 15428
rect 11256 15416 11284 15447
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 11698 15484 11704 15496
rect 11659 15456 11704 15484
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15484 11943 15487
rect 12452 15484 12480 15524
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 13096 15552 13124 15592
rect 13096 15524 13216 15552
rect 11931 15456 12480 15484
rect 12529 15487 12587 15493
rect 11931 15453 11943 15456
rect 11885 15447 11943 15453
rect 12529 15453 12541 15487
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 12544 15416 12572 15447
rect 12986 15444 12992 15496
rect 13044 15484 13050 15496
rect 13188 15493 13216 15524
rect 13173 15487 13231 15493
rect 13044 15456 13089 15484
rect 13044 15444 13050 15456
rect 13173 15453 13185 15487
rect 13219 15453 13231 15487
rect 13173 15447 13231 15453
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15453 14427 15487
rect 14369 15447 14427 15453
rect 15565 15487 15623 15493
rect 15565 15453 15577 15487
rect 15611 15484 15623 15487
rect 15838 15484 15844 15496
rect 15611 15456 15844 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 13354 15416 13360 15428
rect 10652 15388 11284 15416
rect 11348 15388 12112 15416
rect 12544 15388 13360 15416
rect 10652 15376 10658 15388
rect 11348 15348 11376 15388
rect 10428 15320 11376 15348
rect 11514 15308 11520 15360
rect 11572 15348 11578 15360
rect 11698 15348 11704 15360
rect 11572 15320 11704 15348
rect 11572 15308 11578 15320
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 11793 15351 11851 15357
rect 11793 15317 11805 15351
rect 11839 15348 11851 15351
rect 11974 15348 11980 15360
rect 11839 15320 11980 15348
rect 11839 15317 11851 15320
rect 11793 15311 11851 15317
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12084 15348 12112 15388
rect 13354 15376 13360 15388
rect 13412 15376 13418 15428
rect 14384 15348 14412 15447
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 12084 15320 14412 15348
rect 15749 15351 15807 15357
rect 15749 15317 15761 15351
rect 15795 15348 15807 15351
rect 16666 15348 16672 15360
rect 15795 15320 16672 15348
rect 15795 15317 15807 15320
rect 15749 15311 15807 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 1104 15258 16836 15280
rect 1104 15206 4898 15258
rect 4950 15206 4962 15258
rect 5014 15206 5026 15258
rect 5078 15206 5090 15258
rect 5142 15206 5154 15258
rect 5206 15206 8846 15258
rect 8898 15206 8910 15258
rect 8962 15206 8974 15258
rect 9026 15206 9038 15258
rect 9090 15206 9102 15258
rect 9154 15206 12794 15258
rect 12846 15206 12858 15258
rect 12910 15206 12922 15258
rect 12974 15206 12986 15258
rect 13038 15206 13050 15258
rect 13102 15206 16836 15258
rect 1104 15184 16836 15206
rect 1397 15147 1455 15153
rect 1397 15113 1409 15147
rect 1443 15144 1455 15147
rect 1854 15144 1860 15156
rect 1443 15116 1860 15144
rect 1443 15113 1455 15116
rect 1397 15107 1455 15113
rect 1854 15104 1860 15116
rect 1912 15104 1918 15156
rect 2222 15104 2228 15156
rect 2280 15144 2286 15156
rect 4522 15144 4528 15156
rect 2280 15116 4528 15144
rect 2280 15104 2286 15116
rect 4522 15104 4528 15116
rect 4580 15104 4586 15156
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 5408 15116 7052 15144
rect 5408 15104 5414 15116
rect 2682 15076 2688 15088
rect 1688 15048 2688 15076
rect 1578 15008 1584 15020
rect 1636 15017 1642 15020
rect 1500 14980 1584 15008
rect 1578 14968 1584 14980
rect 1636 15008 1648 15017
rect 1688 15008 1716 15048
rect 2682 15036 2688 15048
rect 2740 15036 2746 15088
rect 2958 15036 2964 15088
rect 3016 15076 3022 15088
rect 4614 15076 4620 15088
rect 3016 15048 4620 15076
rect 3016 15036 3022 15048
rect 4614 15036 4620 15048
rect 4672 15085 4678 15088
rect 4672 15079 4736 15085
rect 4672 15045 4690 15079
rect 4724 15076 4736 15079
rect 5902 15076 5908 15088
rect 4724 15048 5908 15076
rect 4724 15045 4736 15048
rect 4672 15039 4736 15045
rect 4672 15036 4678 15039
rect 5902 15036 5908 15048
rect 5960 15036 5966 15088
rect 6270 15036 6276 15088
rect 6328 15076 6334 15088
rect 6917 15079 6975 15085
rect 6917 15076 6929 15079
rect 6328 15048 6929 15076
rect 6328 15036 6334 15048
rect 6917 15045 6929 15048
rect 6963 15045 6975 15079
rect 7024 15076 7052 15116
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 9030 15144 9036 15156
rect 8352 15116 9036 15144
rect 8352 15104 8358 15116
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9306 15104 9312 15156
rect 9364 15144 9370 15156
rect 11330 15144 11336 15156
rect 9364 15116 11336 15144
rect 9364 15104 9370 15116
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 11698 15144 11704 15156
rect 11659 15116 11704 15144
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 13538 15144 13544 15156
rect 12308 15116 13544 15144
rect 12308 15104 12314 15116
rect 13538 15104 13544 15116
rect 13596 15104 13602 15156
rect 13722 15104 13728 15156
rect 13780 15144 13786 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 13780 15116 13829 15144
rect 13780 15104 13786 15116
rect 13817 15113 13829 15116
rect 13863 15113 13875 15147
rect 15654 15144 15660 15156
rect 15615 15116 15660 15144
rect 13817 15107 13875 15113
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 8021 15079 8079 15085
rect 8021 15076 8033 15079
rect 7024 15048 8033 15076
rect 6917 15039 6975 15045
rect 8021 15045 8033 15048
rect 8067 15045 8079 15079
rect 8021 15039 8079 15045
rect 8110 15036 8116 15088
rect 8168 15076 8174 15088
rect 10413 15079 10471 15085
rect 10413 15076 10425 15079
rect 8168 15048 10425 15076
rect 8168 15036 8174 15048
rect 10413 15045 10425 15048
rect 10459 15045 10471 15079
rect 10413 15039 10471 15045
rect 10520 15048 11376 15076
rect 10520 15020 10548 15048
rect 1854 15008 1860 15020
rect 1636 14980 1716 15008
rect 1815 14980 1860 15008
rect 1636 14971 1648 14980
rect 1636 14968 1642 14971
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 2314 15008 2320 15020
rect 2087 14980 2320 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 2866 15017 2872 15020
rect 2860 15008 2872 15017
rect 2424 14980 2872 15008
rect 1762 14900 1768 14952
rect 1820 14940 1826 14952
rect 2424 14940 2452 14980
rect 2860 14971 2872 14980
rect 2866 14968 2872 14971
rect 2924 14968 2930 15020
rect 6457 15011 6515 15017
rect 6457 14977 6469 15011
rect 6503 15008 6515 15011
rect 6546 15008 6552 15020
rect 6503 14980 6552 15008
rect 6503 14977 6515 14980
rect 6457 14971 6515 14977
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 6638 14968 6644 15020
rect 6696 15008 6702 15020
rect 7190 15008 7196 15020
rect 6696 14980 6741 15008
rect 7151 14980 7196 15008
rect 6696 14968 6702 14980
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 8294 14968 8300 15020
rect 8352 15008 8358 15020
rect 9306 15008 9312 15020
rect 8352 14980 9312 15008
rect 8352 14968 8358 14980
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 10229 15011 10287 15017
rect 9732 14980 10180 15008
rect 9732 14968 9738 14980
rect 1820 14912 2452 14940
rect 1820 14900 1826 14912
rect 2590 14900 2596 14952
rect 2648 14940 2654 14952
rect 2648 14912 2693 14940
rect 2648 14900 2654 14912
rect 4154 14900 4160 14952
rect 4212 14940 4218 14952
rect 4433 14943 4491 14949
rect 4433 14940 4445 14943
rect 4212 14912 4445 14940
rect 4212 14900 4218 14912
rect 4433 14909 4445 14912
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 6178 14900 6184 14952
rect 6236 14940 6242 14952
rect 6656 14940 6684 14968
rect 6236 14912 6684 14940
rect 6236 14900 6242 14912
rect 7466 14900 7472 14952
rect 7524 14940 7530 14952
rect 9950 14940 9956 14952
rect 7524 14912 9956 14940
rect 7524 14900 7530 14912
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 10152 14940 10180 14980
rect 10229 14977 10241 15011
rect 10275 15008 10287 15011
rect 10318 15008 10324 15020
rect 10275 14980 10324 15008
rect 10275 14977 10287 14980
rect 10229 14971 10287 14977
rect 10318 14968 10324 14980
rect 10376 14968 10382 15020
rect 10502 15008 10508 15020
rect 10463 14980 10508 15008
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 14977 10655 15011
rect 11348 15008 11376 15048
rect 11422 15036 11428 15088
rect 11480 15076 11486 15088
rect 11517 15079 11575 15085
rect 11517 15076 11529 15079
rect 11480 15048 11529 15076
rect 11480 15036 11486 15048
rect 11517 15045 11529 15048
rect 11563 15045 11575 15079
rect 15930 15076 15936 15088
rect 11517 15039 11575 15045
rect 11992 15048 15936 15076
rect 11992 15017 12020 15048
rect 15930 15036 15936 15048
rect 15988 15036 15994 15088
rect 12434 15017 12440 15020
rect 11977 15011 12035 15017
rect 11348 14980 11928 15008
rect 10597 14971 10655 14977
rect 10612 14940 10640 14971
rect 11698 14940 11704 14952
rect 10152 14912 11704 14940
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 11900 14940 11928 14980
rect 11977 14977 11989 15011
rect 12023 14977 12035 15011
rect 11977 14971 12035 14977
rect 12429 14971 12440 15017
rect 12492 15008 12498 15020
rect 12492 14980 12529 15008
rect 12434 14968 12440 14971
rect 12492 14968 12498 14980
rect 12894 14968 12900 15020
rect 12952 15008 12958 15020
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 12952 14980 13093 15008
rect 12952 14968 12958 14980
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13722 15008 13728 15020
rect 13683 14980 13728 15008
rect 13081 14971 13139 14977
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 14921 15011 14979 15017
rect 14921 15008 14933 15011
rect 13872 14980 14933 15008
rect 13872 14968 13878 14980
rect 14921 14977 14933 14980
rect 14967 14977 14979 15011
rect 15562 15008 15568 15020
rect 15523 14980 15568 15008
rect 14921 14971 14979 14977
rect 15562 14968 15568 14980
rect 15620 14968 15626 15020
rect 14182 14940 14188 14952
rect 11900 14912 14188 14940
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 1578 14832 1584 14884
rect 1636 14872 1642 14884
rect 2608 14872 2636 14900
rect 1636 14844 2636 14872
rect 1636 14832 1642 14844
rect 5626 14832 5632 14884
rect 5684 14872 5690 14884
rect 10594 14872 10600 14884
rect 5684 14844 10600 14872
rect 5684 14832 5690 14844
rect 10594 14832 10600 14844
rect 10652 14832 10658 14884
rect 12621 14875 12679 14881
rect 12621 14872 12633 14875
rect 10704 14844 12633 14872
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 3973 14807 4031 14813
rect 3973 14804 3985 14807
rect 1820 14776 3985 14804
rect 1820 14764 1826 14776
rect 3973 14773 3985 14776
rect 4019 14773 4031 14807
rect 3973 14767 4031 14773
rect 4154 14764 4160 14816
rect 4212 14804 4218 14816
rect 5813 14807 5871 14813
rect 5813 14804 5825 14807
rect 4212 14776 5825 14804
rect 4212 14764 4218 14776
rect 5813 14773 5825 14776
rect 5859 14773 5871 14807
rect 5813 14767 5871 14773
rect 5902 14764 5908 14816
rect 5960 14804 5966 14816
rect 8846 14804 8852 14816
rect 5960 14776 8852 14804
rect 5960 14764 5966 14776
rect 8846 14764 8852 14776
rect 8904 14764 8910 14816
rect 8938 14764 8944 14816
rect 8996 14804 9002 14816
rect 9309 14807 9367 14813
rect 9309 14804 9321 14807
rect 8996 14776 9321 14804
rect 8996 14764 9002 14776
rect 9309 14773 9321 14776
rect 9355 14773 9367 14807
rect 9309 14767 9367 14773
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 10704 14804 10732 14844
rect 12621 14841 12633 14844
rect 12667 14841 12679 14875
rect 12621 14835 12679 14841
rect 15105 14875 15163 14881
rect 15105 14841 15117 14875
rect 15151 14872 15163 14875
rect 15654 14872 15660 14884
rect 15151 14844 15660 14872
rect 15151 14841 15163 14844
rect 15105 14835 15163 14841
rect 15654 14832 15660 14844
rect 15712 14832 15718 14884
rect 9732 14776 10732 14804
rect 10781 14807 10839 14813
rect 9732 14764 9738 14776
rect 10781 14773 10793 14807
rect 10827 14804 10839 14807
rect 11606 14804 11612 14816
rect 10827 14776 11612 14804
rect 10827 14773 10839 14776
rect 10781 14767 10839 14773
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 11701 14807 11759 14813
rect 11701 14773 11713 14807
rect 11747 14804 11759 14807
rect 12434 14804 12440 14816
rect 11747 14776 12440 14804
rect 11747 14773 11759 14776
rect 11701 14767 11759 14773
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 13262 14804 13268 14816
rect 13223 14776 13268 14804
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 1104 14714 16836 14736
rect 1104 14662 2924 14714
rect 2976 14662 2988 14714
rect 3040 14662 3052 14714
rect 3104 14662 3116 14714
rect 3168 14662 3180 14714
rect 3232 14662 6872 14714
rect 6924 14662 6936 14714
rect 6988 14662 7000 14714
rect 7052 14662 7064 14714
rect 7116 14662 7128 14714
rect 7180 14662 10820 14714
rect 10872 14662 10884 14714
rect 10936 14662 10948 14714
rect 11000 14662 11012 14714
rect 11064 14662 11076 14714
rect 11128 14662 14768 14714
rect 14820 14662 14832 14714
rect 14884 14662 14896 14714
rect 14948 14662 14960 14714
rect 15012 14662 15024 14714
rect 15076 14662 16836 14714
rect 1104 14640 16836 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 3237 14603 3295 14609
rect 3237 14600 3249 14603
rect 1912 14572 3249 14600
rect 1912 14560 1918 14572
rect 3237 14569 3249 14572
rect 3283 14569 3295 14603
rect 7006 14600 7012 14612
rect 3237 14563 3295 14569
rect 4264 14572 7012 14600
rect 1578 14424 1584 14476
rect 1636 14464 1642 14476
rect 4264 14473 4292 14572
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 7282 14600 7288 14612
rect 7156 14572 7288 14600
rect 7156 14560 7162 14572
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 7469 14603 7527 14609
rect 7469 14569 7481 14603
rect 7515 14600 7527 14603
rect 7742 14600 7748 14612
rect 7515 14572 7748 14600
rect 7515 14569 7527 14572
rect 7469 14563 7527 14569
rect 5626 14532 5632 14544
rect 5587 14504 5632 14532
rect 5626 14492 5632 14504
rect 5684 14492 5690 14544
rect 1857 14467 1915 14473
rect 1857 14464 1869 14467
rect 1636 14436 1869 14464
rect 1636 14424 1642 14436
rect 1857 14433 1869 14436
rect 1903 14433 1915 14467
rect 1857 14427 1915 14433
rect 4249 14467 4307 14473
rect 4249 14433 4261 14467
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 4516 14399 4574 14405
rect 4516 14365 4528 14399
rect 4562 14396 4574 14399
rect 5902 14396 5908 14408
rect 4562 14368 5908 14396
rect 4562 14365 4574 14368
rect 4516 14359 4574 14365
rect 5902 14356 5908 14368
rect 5960 14356 5966 14408
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14396 6147 14399
rect 6135 14368 6592 14396
rect 6135 14365 6147 14368
rect 6089 14359 6147 14365
rect 6564 14340 6592 14368
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 7484 14396 7512 14563
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 11425 14603 11483 14609
rect 11425 14600 11437 14603
rect 8904 14572 11437 14600
rect 8904 14560 8910 14572
rect 11425 14569 11437 14572
rect 11471 14569 11483 14603
rect 11425 14563 11483 14569
rect 11514 14560 11520 14612
rect 11572 14600 11578 14612
rect 11572 14572 11928 14600
rect 11572 14560 11578 14572
rect 7432 14368 7512 14396
rect 7760 14504 8708 14532
rect 7432 14356 7438 14368
rect 1394 14288 1400 14340
rect 1452 14328 1458 14340
rect 1578 14328 1584 14340
rect 1452 14300 1584 14328
rect 1452 14288 1458 14300
rect 1578 14288 1584 14300
rect 1636 14328 1642 14340
rect 2102 14331 2160 14337
rect 2102 14328 2114 14331
rect 1636 14300 2114 14328
rect 1636 14288 1642 14300
rect 2102 14297 2114 14300
rect 2148 14297 2160 14331
rect 2102 14291 2160 14297
rect 6356 14331 6414 14337
rect 6356 14297 6368 14331
rect 6402 14328 6414 14331
rect 6454 14328 6460 14340
rect 6402 14300 6460 14328
rect 6402 14297 6414 14300
rect 6356 14291 6414 14297
rect 6454 14288 6460 14300
rect 6512 14288 6518 14340
rect 6546 14288 6552 14340
rect 6604 14288 6610 14340
rect 7760 14328 7788 14504
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 8570 14464 8576 14476
rect 8352 14436 8576 14464
rect 8352 14424 8358 14436
rect 8570 14424 8576 14436
rect 8628 14424 8634 14476
rect 8680 14464 8708 14504
rect 8754 14492 8760 14544
rect 8812 14532 8818 14544
rect 9030 14532 9036 14544
rect 8812 14504 9036 14532
rect 8812 14492 8818 14504
rect 9030 14492 9036 14504
rect 9088 14492 9094 14544
rect 9122 14492 9128 14544
rect 9180 14532 9186 14544
rect 10229 14535 10287 14541
rect 9180 14504 9260 14532
rect 9180 14492 9186 14504
rect 9232 14473 9260 14504
rect 10229 14501 10241 14535
rect 10275 14532 10287 14535
rect 10410 14532 10416 14544
rect 10275 14504 10416 14532
rect 10275 14501 10287 14504
rect 10229 14495 10287 14501
rect 10410 14492 10416 14504
rect 10468 14492 10474 14544
rect 10594 14492 10600 14544
rect 10652 14532 10658 14544
rect 11900 14532 11928 14572
rect 12066 14560 12072 14612
rect 12124 14600 12130 14612
rect 12529 14603 12587 14609
rect 12529 14600 12541 14603
rect 12124 14572 12541 14600
rect 12124 14560 12130 14572
rect 12529 14569 12541 14572
rect 12575 14569 12587 14603
rect 12529 14563 12587 14569
rect 12713 14603 12771 14609
rect 12713 14569 12725 14603
rect 12759 14600 12771 14603
rect 12894 14600 12900 14612
rect 12759 14572 12900 14600
rect 12759 14569 12771 14572
rect 12713 14563 12771 14569
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 14737 14603 14795 14609
rect 14737 14600 14749 14603
rect 14332 14572 14749 14600
rect 14332 14560 14338 14572
rect 14737 14569 14749 14572
rect 14783 14569 14795 14603
rect 14737 14563 14795 14569
rect 10652 14504 11836 14532
rect 11900 14504 15608 14532
rect 10652 14492 10658 14504
rect 9217 14467 9275 14473
rect 8680 14436 9168 14464
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14396 8079 14399
rect 8478 14396 8484 14408
rect 8067 14368 8484 14396
rect 8067 14365 8079 14368
rect 8021 14359 8079 14365
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 8941 14399 8999 14405
rect 8941 14365 8953 14399
rect 8987 14396 8999 14399
rect 9030 14396 9036 14408
rect 8987 14368 9036 14396
rect 8987 14365 8999 14368
rect 8941 14359 8999 14365
rect 9030 14356 9036 14368
rect 9088 14356 9094 14408
rect 9140 14396 9168 14436
rect 9217 14433 9229 14467
rect 9263 14433 9275 14467
rect 9217 14427 9275 14433
rect 9858 14424 9864 14476
rect 9916 14464 9922 14476
rect 9916 14436 10824 14464
rect 9916 14424 9922 14436
rect 10689 14399 10747 14405
rect 9140 14390 10640 14396
rect 10689 14390 10701 14399
rect 9140 14368 10701 14390
rect 10612 14365 10701 14368
rect 10735 14365 10747 14399
rect 10796 14396 10824 14436
rect 10870 14424 10876 14476
rect 10928 14464 10934 14476
rect 11808 14464 11836 14504
rect 12526 14464 12532 14476
rect 10928 14436 10973 14464
rect 11440 14436 11740 14464
rect 10928 14424 10934 14436
rect 11440 14408 11468 14436
rect 11422 14396 11428 14408
rect 10796 14368 11428 14396
rect 10612 14362 10747 14365
rect 10689 14359 10747 14362
rect 11422 14356 11428 14368
rect 11480 14356 11486 14408
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 6656 14300 7788 14328
rect 8205 14331 8263 14337
rect 1210 14220 1216 14272
rect 1268 14260 1274 14272
rect 1854 14260 1860 14272
rect 1268 14232 1860 14260
rect 1268 14220 1274 14232
rect 1854 14220 1860 14232
rect 1912 14220 1918 14272
rect 2406 14220 2412 14272
rect 2464 14260 2470 14272
rect 6656 14260 6684 14300
rect 8205 14297 8217 14331
rect 8251 14328 8263 14331
rect 8570 14328 8576 14340
rect 8251 14300 8576 14328
rect 8251 14297 8263 14300
rect 8205 14291 8263 14297
rect 8570 14288 8576 14300
rect 8628 14288 8634 14340
rect 8662 14288 8668 14340
rect 8720 14328 8726 14340
rect 9214 14328 9220 14340
rect 8720 14300 9220 14328
rect 8720 14288 8726 14300
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 9766 14288 9772 14340
rect 9824 14328 9830 14340
rect 9824 14300 10732 14328
rect 9824 14288 9830 14300
rect 10704 14272 10732 14300
rect 11238 14288 11244 14340
rect 11296 14328 11302 14340
rect 11514 14328 11520 14340
rect 11296 14300 11520 14328
rect 11296 14288 11302 14300
rect 11514 14288 11520 14300
rect 11572 14328 11578 14340
rect 11624 14328 11652 14359
rect 11572 14300 11652 14328
rect 11712 14328 11740 14436
rect 11808 14436 12532 14464
rect 11808 14405 11836 14436
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 13357 14467 13415 14473
rect 13357 14464 13369 14467
rect 12768 14436 13369 14464
rect 12768 14424 12774 14436
rect 13357 14433 13369 14436
rect 13403 14433 13415 14467
rect 13357 14427 13415 14433
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 13596 14436 15424 14464
rect 13596 14424 13602 14436
rect 11793 14399 11851 14405
rect 11793 14365 11805 14399
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14396 11943 14399
rect 12158 14396 12164 14408
rect 11931 14368 12164 14396
rect 11931 14365 11943 14368
rect 11885 14359 11943 14365
rect 12158 14356 12164 14368
rect 12216 14396 12222 14408
rect 12216 14368 12472 14396
rect 12216 14356 12222 14368
rect 12345 14331 12403 14337
rect 12345 14328 12357 14331
rect 11712 14300 12357 14328
rect 11572 14288 11578 14300
rect 12345 14297 12357 14300
rect 12391 14297 12403 14331
rect 12444 14328 12472 14368
rect 13170 14356 13176 14408
rect 13228 14396 13234 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 13228 14368 13277 14396
rect 13228 14356 13234 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 13446 14396 13452 14408
rect 13407 14368 13452 14396
rect 13265 14359 13323 14365
rect 13446 14356 13452 14368
rect 13504 14396 13510 14408
rect 13630 14396 13636 14408
rect 13504 14368 13636 14396
rect 13504 14356 13510 14368
rect 13630 14356 13636 14368
rect 13688 14356 13694 14408
rect 13998 14356 14004 14408
rect 14056 14396 14062 14408
rect 14277 14399 14335 14405
rect 14277 14396 14289 14399
rect 14056 14368 14289 14396
rect 14056 14356 14062 14368
rect 14277 14365 14289 14368
rect 14323 14365 14335 14399
rect 14918 14396 14924 14408
rect 14879 14368 14924 14396
rect 14277 14359 14335 14365
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 15396 14405 15424 14436
rect 15580 14405 15608 14504
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14365 15439 14399
rect 15381 14359 15439 14365
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 14642 14328 14648 14340
rect 12444 14300 14648 14328
rect 12345 14291 12403 14297
rect 14642 14288 14648 14300
rect 14700 14288 14706 14340
rect 2464 14232 6684 14260
rect 2464 14220 2470 14232
rect 7190 14220 7196 14272
rect 7248 14260 7254 14272
rect 9398 14260 9404 14272
rect 7248 14232 9404 14260
rect 7248 14220 7254 14232
rect 9398 14220 9404 14232
rect 9456 14220 9462 14272
rect 9490 14220 9496 14272
rect 9548 14260 9554 14272
rect 10597 14263 10655 14269
rect 10597 14260 10609 14263
rect 9548 14232 10609 14260
rect 9548 14220 9554 14232
rect 10597 14229 10609 14232
rect 10643 14229 10655 14263
rect 10597 14223 10655 14229
rect 10686 14220 10692 14272
rect 10744 14220 10750 14272
rect 11330 14220 11336 14272
rect 11388 14260 11394 14272
rect 11606 14260 11612 14272
rect 11388 14232 11612 14260
rect 11388 14220 11394 14232
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 11698 14220 11704 14272
rect 11756 14260 11762 14272
rect 12529 14263 12587 14269
rect 12529 14260 12541 14263
rect 11756 14232 12541 14260
rect 11756 14220 11762 14232
rect 12529 14229 12541 14232
rect 12575 14260 12587 14263
rect 13630 14260 13636 14272
rect 12575 14232 13636 14260
rect 12575 14229 12587 14232
rect 12529 14223 12587 14229
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14093 14263 14151 14269
rect 14093 14260 14105 14263
rect 13872 14232 14105 14260
rect 13872 14220 13878 14232
rect 14093 14229 14105 14232
rect 14139 14229 14151 14263
rect 14093 14223 14151 14229
rect 15010 14220 15016 14272
rect 15068 14260 15074 14272
rect 15473 14263 15531 14269
rect 15473 14260 15485 14263
rect 15068 14232 15485 14260
rect 15068 14220 15074 14232
rect 15473 14229 15485 14232
rect 15519 14229 15531 14263
rect 15473 14223 15531 14229
rect 1104 14170 16836 14192
rect 1104 14118 4898 14170
rect 4950 14118 4962 14170
rect 5014 14118 5026 14170
rect 5078 14118 5090 14170
rect 5142 14118 5154 14170
rect 5206 14118 8846 14170
rect 8898 14118 8910 14170
rect 8962 14118 8974 14170
rect 9026 14118 9038 14170
rect 9090 14118 9102 14170
rect 9154 14118 12794 14170
rect 12846 14118 12858 14170
rect 12910 14118 12922 14170
rect 12974 14118 12986 14170
rect 13038 14118 13050 14170
rect 13102 14118 16836 14170
rect 1104 14096 16836 14118
rect 1210 14016 1216 14068
rect 1268 14056 1274 14068
rect 5169 14059 5227 14065
rect 1268 14028 5028 14056
rect 1268 14016 1274 14028
rect 1118 13948 1124 14000
rect 1176 13988 1182 14000
rect 1394 13988 1400 14000
rect 1176 13960 1400 13988
rect 1176 13948 1182 13960
rect 1394 13948 1400 13960
rect 1452 13948 1458 14000
rect 1762 13988 1768 14000
rect 1723 13960 1768 13988
rect 1762 13948 1768 13960
rect 1820 13948 1826 14000
rect 1857 13991 1915 13997
rect 1857 13957 1869 13991
rect 1903 13988 1915 13991
rect 2222 13988 2228 14000
rect 1903 13960 2228 13988
rect 1903 13957 1915 13960
rect 1857 13951 1915 13957
rect 2222 13948 2228 13960
rect 2280 13948 2286 14000
rect 750 13880 756 13932
rect 808 13880 814 13932
rect 2406 13920 2412 13932
rect 1964 13892 2412 13920
rect 768 13852 796 13880
rect 1762 13852 1768 13864
rect 768 13824 1768 13852
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 1397 13787 1455 13793
rect 1397 13753 1409 13787
rect 1443 13784 1455 13787
rect 1964 13784 1992 13892
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 2590 13920 2596 13932
rect 2551 13892 2596 13920
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 3970 13880 3976 13932
rect 4028 13880 4034 13932
rect 5000 13929 5028 14028
rect 5169 14025 5181 14059
rect 5215 14056 5227 14059
rect 6638 14056 6644 14068
rect 5215 14028 6644 14056
rect 5215 14025 5227 14028
rect 5169 14019 5227 14025
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 7558 14016 7564 14068
rect 7616 14056 7622 14068
rect 8938 14056 8944 14068
rect 7616 14028 8944 14056
rect 7616 14016 7622 14028
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9950 14056 9956 14068
rect 9048 14028 9956 14056
rect 7285 13991 7343 13997
rect 7285 13957 7297 13991
rect 7331 13988 7343 13991
rect 7466 13988 7472 14000
rect 7331 13960 7472 13988
rect 7331 13957 7343 13960
rect 7285 13951 7343 13957
rect 7466 13948 7472 13960
rect 7524 13948 7530 14000
rect 7742 13948 7748 14000
rect 7800 13988 7806 14000
rect 9048 13988 9076 14028
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10275 14059 10333 14065
rect 10275 14025 10287 14059
rect 10321 14025 10333 14059
rect 10275 14019 10333 14025
rect 7800 13960 9076 13988
rect 7800 13948 7806 13960
rect 9122 13948 9128 14000
rect 9180 13988 9186 14000
rect 10290 13988 10318 14019
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 11112 14028 12909 14056
rect 11112 14016 11118 14028
rect 12897 14025 12909 14028
rect 12943 14025 12955 14059
rect 12897 14019 12955 14025
rect 13998 14016 14004 14068
rect 14056 14056 14062 14068
rect 14056 14028 14780 14056
rect 14056 14016 14062 14028
rect 9180 13960 10318 13988
rect 9180 13948 9186 13960
rect 10502 13948 10508 14000
rect 10560 13988 10566 14000
rect 10560 13960 12020 13988
rect 10560 13948 10566 13960
rect 4985 13923 5043 13929
rect 4985 13889 4997 13923
rect 5031 13889 5043 13923
rect 4985 13883 5043 13889
rect 5629 13923 5687 13929
rect 5629 13889 5641 13923
rect 5675 13889 5687 13923
rect 5810 13920 5816 13932
rect 5771 13892 5816 13920
rect 5629 13883 5687 13889
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 1443 13756 1992 13784
rect 2056 13784 2084 13815
rect 2406 13784 2412 13796
rect 2056 13756 2412 13784
rect 1443 13753 1455 13756
rect 1397 13747 1455 13753
rect 2406 13744 2412 13756
rect 2464 13744 2470 13796
rect 1486 13676 1492 13728
rect 1544 13716 1550 13728
rect 2222 13716 2228 13728
rect 1544 13688 2228 13716
rect 1544 13676 1550 13688
rect 2222 13676 2228 13688
rect 2280 13716 2286 13728
rect 2608 13716 2636 13880
rect 2958 13812 2964 13864
rect 3016 13852 3022 13864
rect 5644 13852 5672 13883
rect 5810 13880 5816 13892
rect 5868 13880 5874 13932
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 7098 13920 7104 13932
rect 6512 13892 7104 13920
rect 6512 13880 6518 13892
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 7248 13892 7389 13920
rect 7248 13880 7254 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 9398 13920 9404 13932
rect 7883 13892 9404 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 10226 13880 10232 13932
rect 10284 13920 10290 13932
rect 11992 13929 12020 13960
rect 12066 13948 12072 14000
rect 12124 13988 12130 14000
rect 13906 13988 13912 14000
rect 12124 13960 12572 13988
rect 12124 13948 12130 13960
rect 12544 13929 12572 13960
rect 13740 13960 13912 13988
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 10284 13892 11529 13920
rect 10284 13880 10290 13892
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12529 13923 12587 13929
rect 12529 13889 12541 13923
rect 12575 13889 12587 13923
rect 12710 13920 12716 13932
rect 12671 13892 12716 13920
rect 12529 13883 12587 13889
rect 3016 13824 5672 13852
rect 6917 13855 6975 13861
rect 3016 13812 3022 13824
rect 6917 13821 6929 13855
rect 6963 13852 6975 13855
rect 9490 13852 9496 13864
rect 6963 13824 9496 13852
rect 6963 13821 6975 13824
rect 6917 13815 6975 13821
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 9858 13852 9864 13864
rect 9692 13824 9864 13852
rect 4341 13787 4399 13793
rect 4341 13753 4353 13787
rect 4387 13753 4399 13787
rect 4341 13747 4399 13753
rect 2866 13725 2872 13728
rect 2856 13719 2872 13725
rect 2856 13716 2868 13719
rect 2280 13688 2636 13716
rect 2779 13688 2868 13716
rect 2280 13676 2286 13688
rect 2856 13685 2868 13688
rect 2924 13716 2930 13728
rect 3970 13716 3976 13728
rect 2924 13688 3976 13716
rect 2856 13679 2872 13685
rect 2866 13676 2872 13679
rect 2924 13676 2930 13688
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4356 13716 4384 13747
rect 7006 13744 7012 13796
rect 7064 13784 7070 13796
rect 7064 13756 7880 13784
rect 7064 13744 7070 13756
rect 4706 13716 4712 13728
rect 4356 13688 4712 13716
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 5629 13719 5687 13725
rect 5629 13685 5641 13719
rect 5675 13716 5687 13719
rect 7190 13716 7196 13728
rect 5675 13688 7196 13716
rect 5675 13685 5687 13688
rect 5629 13679 5687 13685
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 7852 13716 7880 13756
rect 8662 13744 8668 13796
rect 8720 13784 8726 13796
rect 9692 13784 9720 13824
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 9950 13812 9956 13864
rect 10008 13852 10014 13864
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 10008 13824 10057 13852
rect 10008 13812 10014 13824
rect 10045 13821 10057 13824
rect 10091 13852 10103 13855
rect 10410 13852 10416 13864
rect 10091 13824 10416 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10410 13812 10416 13824
rect 10468 13812 10474 13864
rect 11072 13824 11284 13852
rect 8720 13756 9720 13784
rect 8720 13744 8726 13756
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 11072 13784 11100 13824
rect 9824 13756 11100 13784
rect 11256 13784 11284 13824
rect 11330 13812 11336 13864
rect 11388 13852 11394 13864
rect 11716 13852 11744 13883
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12952 13892 13001 13920
rect 12952 13880 12958 13892
rect 12989 13889 13001 13892
rect 13035 13920 13047 13923
rect 13078 13920 13084 13932
rect 13035 13892 13084 13920
rect 13035 13889 13047 13892
rect 12989 13883 13047 13889
rect 13078 13880 13084 13892
rect 13136 13880 13142 13932
rect 13740 13929 13768 13960
rect 13906 13948 13912 13960
rect 13964 13988 13970 14000
rect 14458 13988 14464 14000
rect 13964 13960 14464 13988
rect 13964 13948 13970 13960
rect 14458 13948 14464 13960
rect 14516 13988 14522 14000
rect 14752 13997 14780 14028
rect 14737 13991 14795 13997
rect 14516 13960 14596 13988
rect 14516 13948 14522 13960
rect 14568 13929 14596 13960
rect 14737 13957 14749 13991
rect 14783 13957 14795 13991
rect 14737 13951 14795 13957
rect 15194 13948 15200 14000
rect 15252 13988 15258 14000
rect 15657 13991 15715 13997
rect 15657 13988 15669 13991
rect 15252 13960 15669 13988
rect 15252 13948 15258 13960
rect 15657 13957 15669 13960
rect 15703 13957 15715 13991
rect 15657 13951 15715 13957
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 14369 13923 14427 13929
rect 14369 13920 14381 13923
rect 13725 13883 13783 13889
rect 13832 13892 14381 13920
rect 11388 13824 11744 13852
rect 11885 13855 11943 13861
rect 11388 13812 11394 13824
rect 11885 13821 11897 13855
rect 11931 13852 11943 13855
rect 12066 13852 12072 13864
rect 11931 13824 12072 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 13556 13852 13584 13883
rect 13832 13852 13860 13892
rect 14369 13889 14381 13892
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 12860 13824 13860 13852
rect 13909 13855 13967 13861
rect 12860 13812 12866 13824
rect 13909 13821 13921 13855
rect 13955 13852 13967 13855
rect 13998 13852 14004 13864
rect 13955 13824 14004 13852
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 11698 13784 11704 13796
rect 11256 13756 11704 13784
rect 9824 13744 9830 13756
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 11793 13787 11851 13793
rect 11793 13753 11805 13787
rect 11839 13784 11851 13787
rect 14274 13784 14280 13796
rect 11839 13756 14280 13784
rect 11839 13753 11851 13756
rect 11793 13747 11851 13753
rect 14274 13744 14280 13756
rect 14332 13744 14338 13796
rect 15841 13787 15899 13793
rect 15841 13753 15853 13787
rect 15887 13784 15899 13787
rect 16298 13784 16304 13796
rect 15887 13756 16304 13784
rect 15887 13753 15899 13756
rect 15841 13747 15899 13753
rect 16298 13744 16304 13756
rect 16356 13744 16362 13796
rect 8570 13716 8576 13728
rect 7852 13688 8576 13716
rect 8570 13676 8576 13688
rect 8628 13716 8634 13728
rect 9125 13719 9183 13725
rect 9125 13716 9137 13719
rect 8628 13688 9137 13716
rect 8628 13676 8634 13688
rect 9125 13685 9137 13688
rect 9171 13685 9183 13719
rect 9125 13679 9183 13685
rect 9858 13676 9864 13728
rect 9916 13716 9922 13728
rect 10962 13716 10968 13728
rect 9916 13688 10968 13716
rect 9916 13676 9922 13688
rect 10962 13676 10968 13688
rect 11020 13676 11026 13728
rect 11422 13676 11428 13728
rect 11480 13716 11486 13728
rect 12894 13716 12900 13728
rect 11480 13688 12900 13716
rect 11480 13676 11486 13688
rect 12894 13676 12900 13688
rect 12952 13716 12958 13728
rect 16114 13716 16120 13728
rect 12952 13688 16120 13716
rect 12952 13676 12958 13688
rect 16114 13676 16120 13688
rect 16172 13676 16178 13728
rect 1104 13626 16836 13648
rect 1104 13574 2924 13626
rect 2976 13574 2988 13626
rect 3040 13574 3052 13626
rect 3104 13574 3116 13626
rect 3168 13574 3180 13626
rect 3232 13574 6872 13626
rect 6924 13574 6936 13626
rect 6988 13574 7000 13626
rect 7052 13574 7064 13626
rect 7116 13574 7128 13626
rect 7180 13574 10820 13626
rect 10872 13574 10884 13626
rect 10936 13574 10948 13626
rect 11000 13574 11012 13626
rect 11064 13574 11076 13626
rect 11128 13574 14768 13626
rect 14820 13574 14832 13626
rect 14884 13574 14896 13626
rect 14948 13574 14960 13626
rect 15012 13574 15024 13626
rect 15076 13574 16836 13626
rect 1104 13552 16836 13574
rect 1854 13472 1860 13524
rect 1912 13512 1918 13524
rect 3237 13515 3295 13521
rect 3237 13512 3249 13515
rect 1912 13484 3249 13512
rect 1912 13472 1918 13484
rect 3237 13481 3249 13484
rect 3283 13481 3295 13515
rect 5537 13515 5595 13521
rect 3237 13475 3295 13481
rect 3344 13484 5120 13512
rect 2866 13404 2872 13456
rect 2924 13444 2930 13456
rect 3344 13444 3372 13484
rect 2924 13416 3372 13444
rect 2924 13404 2930 13416
rect 3694 13404 3700 13456
rect 3752 13404 3758 13456
rect 5092 13444 5120 13484
rect 5537 13481 5549 13515
rect 5583 13512 5595 13515
rect 5626 13512 5632 13524
rect 5583 13484 5632 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 5626 13472 5632 13484
rect 5684 13512 5690 13524
rect 7006 13512 7012 13524
rect 5684 13484 7012 13512
rect 5684 13472 5690 13484
rect 7006 13472 7012 13484
rect 7064 13472 7070 13524
rect 7282 13472 7288 13524
rect 7340 13512 7346 13524
rect 7558 13512 7564 13524
rect 7340 13484 7564 13512
rect 7340 13472 7346 13484
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 7834 13472 7840 13524
rect 7892 13512 7898 13524
rect 8478 13512 8484 13524
rect 7892 13484 8484 13512
rect 7892 13472 7898 13484
rect 8478 13472 8484 13484
rect 8536 13512 8542 13524
rect 9858 13512 9864 13524
rect 8536 13484 9864 13512
rect 8536 13472 8542 13484
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 11330 13512 11336 13524
rect 10008 13484 11336 13512
rect 10008 13472 10014 13484
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 12069 13515 12127 13521
rect 12069 13481 12081 13515
rect 12115 13512 12127 13515
rect 12158 13512 12164 13524
rect 12115 13484 12164 13512
rect 12115 13481 12127 13484
rect 12069 13475 12127 13481
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 12268 13484 12848 13512
rect 12268 13444 12296 13484
rect 5092 13416 11008 13444
rect 1765 13379 1823 13385
rect 1765 13345 1777 13379
rect 1811 13376 1823 13379
rect 1854 13376 1860 13388
rect 1811 13348 1860 13376
rect 1811 13345 1823 13348
rect 1765 13339 1823 13345
rect 1854 13336 1860 13348
rect 1912 13336 1918 13388
rect 2222 13336 2228 13388
rect 2280 13376 2286 13388
rect 3234 13376 3240 13388
rect 2280 13348 3240 13376
rect 2280 13336 2286 13348
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 1486 13308 1492 13320
rect 1447 13280 1492 13308
rect 1486 13268 1492 13280
rect 1544 13268 1550 13320
rect 3050 13268 3056 13320
rect 3108 13308 3114 13320
rect 3712 13308 3740 13404
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 4522 13376 4528 13388
rect 4111 13348 4528 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 4522 13336 4528 13348
rect 4580 13336 4586 13388
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 5592 13348 6684 13376
rect 5592 13336 5598 13348
rect 3108 13280 3740 13308
rect 3789 13311 3847 13317
rect 3108 13268 3114 13280
rect 3789 13277 3801 13311
rect 3835 13277 3847 13311
rect 5442 13308 5448 13320
rect 5198 13280 5448 13308
rect 3789 13271 3847 13277
rect 2038 13200 2044 13252
rect 2096 13240 2102 13252
rect 2096 13212 2254 13240
rect 2096 13200 2102 13212
rect 3234 13200 3240 13252
rect 3292 13240 3298 13252
rect 3804 13240 3832 13271
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 6656 13317 6684 13348
rect 7282 13336 7288 13388
rect 7340 13376 7346 13388
rect 7834 13376 7840 13388
rect 7340 13348 7840 13376
rect 7340 13336 7346 13348
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 9950 13376 9956 13388
rect 8312 13348 9956 13376
rect 5997 13311 6055 13317
rect 5997 13308 6009 13311
rect 5684 13280 6009 13308
rect 5684 13268 5690 13280
rect 5997 13277 6009 13280
rect 6043 13277 6055 13311
rect 5997 13271 6055 13277
rect 6181 13311 6239 13317
rect 6181 13277 6193 13311
rect 6227 13277 6239 13311
rect 6181 13271 6239 13277
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 3292 13212 3832 13240
rect 6196 13240 6224 13271
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 7466 13308 7472 13320
rect 6788 13280 7472 13308
rect 6788 13268 6794 13280
rect 7466 13268 7472 13280
rect 7524 13268 7530 13320
rect 8202 13240 8208 13252
rect 6196 13212 8208 13240
rect 3292 13200 3298 13212
rect 8202 13200 8208 13212
rect 8260 13240 8266 13252
rect 8312 13240 8340 13348
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10410 13336 10416 13388
rect 10468 13376 10474 13388
rect 10980 13376 11008 13416
rect 11788 13416 12296 13444
rect 11788 13376 11816 13416
rect 12526 13404 12532 13456
rect 12584 13444 12590 13456
rect 12710 13444 12716 13456
rect 12584 13416 12716 13444
rect 12584 13404 12590 13416
rect 12710 13404 12716 13416
rect 12768 13404 12774 13456
rect 12820 13444 12848 13484
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 12952 13484 12997 13512
rect 12952 13472 12958 13484
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 14550 13512 14556 13524
rect 13228 13484 14556 13512
rect 13228 13472 13234 13484
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 14734 13472 14740 13524
rect 14792 13512 14798 13524
rect 15194 13512 15200 13524
rect 14792 13484 15200 13512
rect 14792 13472 14798 13484
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 15657 13515 15715 13521
rect 15657 13512 15669 13515
rect 15436 13484 15669 13512
rect 15436 13472 15442 13484
rect 15657 13481 15669 13484
rect 15703 13481 15715 13515
rect 15657 13475 15715 13481
rect 15013 13447 15071 13453
rect 15013 13444 15025 13447
rect 12820 13416 15025 13444
rect 15013 13413 15025 13416
rect 15059 13413 15071 13447
rect 15013 13407 15071 13413
rect 12434 13376 12440 13388
rect 10468 13348 10916 13376
rect 10980 13348 11816 13376
rect 11900 13348 12440 13376
rect 10468 13336 10474 13348
rect 10888 13320 10916 13348
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 8662 13308 8668 13320
rect 8435 13280 8668 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 8754 13268 8760 13320
rect 8812 13308 8818 13320
rect 9309 13311 9367 13317
rect 9309 13308 9321 13311
rect 8812 13280 9321 13308
rect 8812 13268 8818 13280
rect 9309 13277 9321 13280
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 10870 13268 10876 13320
rect 10928 13268 10934 13320
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 11204 13280 11529 13308
rect 11204 13268 11210 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 11900 13317 11928 13348
rect 12434 13336 12440 13348
rect 12492 13376 12498 13388
rect 12492 13348 12940 13376
rect 12492 13336 12498 13348
rect 11701 13311 11759 13317
rect 11701 13308 11713 13311
rect 11664 13280 11713 13308
rect 11664 13268 11670 13280
rect 11701 13277 11713 13280
rect 11747 13277 11759 13311
rect 11701 13271 11759 13277
rect 11885 13311 11943 13317
rect 11885 13277 11897 13311
rect 11931 13277 11943 13311
rect 12526 13308 12532 13320
rect 12487 13280 12532 13308
rect 11885 13271 11943 13277
rect 12526 13268 12532 13280
rect 12584 13268 12590 13320
rect 8260 13212 8340 13240
rect 8260 13200 8266 13212
rect 8478 13200 8484 13252
rect 8536 13240 8542 13252
rect 8938 13240 8944 13252
rect 8536 13212 8944 13240
rect 8536 13200 8542 13212
rect 8938 13200 8944 13212
rect 8996 13200 9002 13252
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 10778 13240 10784 13252
rect 9088 13212 10784 13240
rect 9088 13200 9094 13212
rect 10778 13200 10784 13212
rect 10836 13200 10842 13252
rect 11057 13243 11115 13249
rect 11057 13209 11069 13243
rect 11103 13209 11115 13243
rect 11057 13203 11115 13209
rect 3050 13132 3056 13184
rect 3108 13172 3114 13184
rect 5442 13172 5448 13184
rect 3108 13144 5448 13172
rect 3108 13132 3114 13144
rect 5442 13132 5448 13144
rect 5500 13172 5506 13184
rect 5902 13172 5908 13184
rect 5500 13144 5908 13172
rect 5500 13132 5506 13144
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 6089 13175 6147 13181
rect 6089 13141 6101 13175
rect 6135 13172 6147 13175
rect 6362 13172 6368 13184
rect 6135 13144 6368 13172
rect 6135 13141 6147 13144
rect 6089 13135 6147 13141
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 7098 13132 7104 13184
rect 7156 13172 7162 13184
rect 9858 13172 9864 13184
rect 7156 13144 9864 13172
rect 7156 13132 7162 13144
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 10410 13132 10416 13184
rect 10468 13172 10474 13184
rect 10962 13172 10968 13184
rect 10468 13144 10968 13172
rect 10468 13132 10474 13144
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 11072 13172 11100 13203
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 12802 13240 12808 13252
rect 11848 13212 11893 13240
rect 11992 13212 12808 13240
rect 11848 13200 11854 13212
rect 11992 13172 12020 13212
rect 12802 13200 12808 13212
rect 12860 13200 12866 13252
rect 12912 13240 12940 13348
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 15749 13379 15807 13385
rect 15749 13376 15761 13379
rect 13044 13348 15761 13376
rect 13044 13336 13050 13348
rect 15749 13345 15761 13348
rect 15795 13345 15807 13379
rect 15749 13339 15807 13345
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13504 13280 14289 13308
rect 13504 13268 13510 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14550 13308 14556 13320
rect 14511 13280 14556 13308
rect 14277 13271 14335 13277
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 15194 13308 15200 13320
rect 15155 13280 15200 13308
rect 15194 13268 15200 13280
rect 15252 13268 15258 13320
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 16022 13308 16028 13320
rect 15703 13280 16028 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 12912 13212 13124 13240
rect 11072 13144 12020 13172
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 13096 13181 13124 13212
rect 13538 13200 13544 13252
rect 13596 13240 13602 13252
rect 14093 13243 14151 13249
rect 14093 13240 14105 13243
rect 13596 13212 14105 13240
rect 13596 13200 13602 13212
rect 14093 13209 14105 13212
rect 14139 13209 14151 13243
rect 14093 13203 14151 13209
rect 12897 13175 12955 13181
rect 12897 13172 12909 13175
rect 12124 13144 12909 13172
rect 12124 13132 12130 13144
rect 12897 13141 12909 13144
rect 12943 13141 12955 13175
rect 12897 13135 12955 13141
rect 13081 13175 13139 13181
rect 13081 13141 13093 13175
rect 13127 13172 13139 13175
rect 13722 13172 13728 13184
rect 13127 13144 13728 13172
rect 13127 13141 13139 13144
rect 13081 13135 13139 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 14182 13132 14188 13184
rect 14240 13172 14246 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 14240 13144 14473 13172
rect 14240 13132 14246 13144
rect 14461 13141 14473 13144
rect 14507 13141 14519 13175
rect 14461 13135 14519 13141
rect 16025 13175 16083 13181
rect 16025 13141 16037 13175
rect 16071 13172 16083 13175
rect 16390 13172 16396 13184
rect 16071 13144 16396 13172
rect 16071 13141 16083 13144
rect 16025 13135 16083 13141
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 1104 13082 16836 13104
rect 1104 13030 4898 13082
rect 4950 13030 4962 13082
rect 5014 13030 5026 13082
rect 5078 13030 5090 13082
rect 5142 13030 5154 13082
rect 5206 13030 8846 13082
rect 8898 13030 8910 13082
rect 8962 13030 8974 13082
rect 9026 13030 9038 13082
rect 9090 13030 9102 13082
rect 9154 13030 12794 13082
rect 12846 13030 12858 13082
rect 12910 13030 12922 13082
rect 12974 13030 12986 13082
rect 13038 13030 13050 13082
rect 13102 13030 16836 13082
rect 1104 13008 16836 13030
rect 474 12928 480 12980
rect 532 12968 538 12980
rect 1118 12968 1124 12980
rect 532 12940 1124 12968
rect 532 12928 538 12940
rect 1118 12928 1124 12940
rect 1176 12928 1182 12980
rect 2130 12928 2136 12980
rect 2188 12928 2194 12980
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 3050 12968 3056 12980
rect 2271 12940 3056 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 4154 12968 4160 12980
rect 3160 12940 4160 12968
rect 2148 12900 2176 12928
rect 2314 12900 2320 12912
rect 2148 12872 2320 12900
rect 2314 12860 2320 12872
rect 2372 12860 2378 12912
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12801 1823 12835
rect 2038 12832 2044 12844
rect 1999 12804 2044 12832
rect 1765 12795 1823 12801
rect 1780 12764 1808 12795
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 2682 12832 2688 12844
rect 2547 12804 2688 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 2961 12835 3019 12841
rect 2961 12801 2973 12835
rect 3007 12832 3019 12835
rect 3160 12832 3188 12940
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4706 12928 4712 12980
rect 4764 12968 4770 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 4764 12940 4813 12968
rect 4764 12928 4770 12940
rect 4801 12937 4813 12940
rect 4847 12937 4859 12971
rect 4801 12931 4859 12937
rect 4890 12928 4896 12980
rect 4948 12968 4954 12980
rect 5350 12968 5356 12980
rect 4948 12940 5356 12968
rect 4948 12928 4954 12940
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 5902 12928 5908 12980
rect 5960 12968 5966 12980
rect 7282 12968 7288 12980
rect 5960 12940 7288 12968
rect 5960 12928 5966 12940
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 7834 12928 7840 12980
rect 7892 12968 7898 12980
rect 9030 12968 9036 12980
rect 7892 12940 9036 12968
rect 7892 12928 7898 12940
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 11517 12971 11575 12977
rect 11517 12968 11529 12971
rect 9180 12940 11529 12968
rect 9180 12928 9186 12940
rect 11517 12937 11529 12940
rect 11563 12937 11575 12971
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11517 12931 11575 12937
rect 11624 12940 11989 12968
rect 5074 12860 5080 12912
rect 5132 12900 5138 12912
rect 5442 12900 5448 12912
rect 5132 12872 5448 12900
rect 5132 12860 5138 12872
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 5537 12903 5595 12909
rect 5537 12869 5549 12903
rect 5583 12900 5595 12903
rect 6178 12900 6184 12912
rect 5583 12872 6184 12900
rect 5583 12869 5595 12872
rect 5537 12863 5595 12869
rect 6178 12860 6184 12872
rect 6236 12860 6242 12912
rect 7558 12900 7564 12912
rect 6288 12872 7564 12900
rect 3007 12804 3188 12832
rect 3007 12801 3019 12804
rect 2961 12795 3019 12801
rect 5166 12792 5172 12844
rect 5224 12832 5230 12844
rect 5261 12835 5319 12841
rect 5261 12832 5273 12835
rect 5224 12804 5273 12832
rect 5224 12792 5230 12804
rect 5261 12801 5273 12804
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12832 5687 12835
rect 5810 12832 5816 12844
rect 5675 12804 5816 12832
rect 5675 12801 5687 12804
rect 5629 12795 5687 12801
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 2222 12764 2228 12776
rect 1780 12736 2228 12764
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 3050 12724 3056 12776
rect 3108 12764 3114 12776
rect 3145 12767 3203 12773
rect 3145 12764 3157 12767
rect 3108 12736 3157 12764
rect 3108 12724 3114 12736
rect 3145 12733 3157 12736
rect 3191 12733 3203 12767
rect 3145 12727 3203 12733
rect 3234 12724 3240 12776
rect 3292 12764 3298 12776
rect 4062 12773 4068 12776
rect 3881 12767 3939 12773
rect 3881 12764 3893 12767
rect 3292 12736 3893 12764
rect 3292 12724 3298 12736
rect 3881 12733 3893 12736
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 4019 12767 4068 12773
rect 4019 12733 4031 12767
rect 4065 12733 4068 12767
rect 4019 12727 4068 12733
rect 4062 12724 4068 12727
rect 4120 12724 4126 12776
rect 4157 12767 4215 12773
rect 4157 12733 4169 12767
rect 4203 12764 4215 12767
rect 4522 12764 4528 12776
rect 4203 12736 4528 12764
rect 4203 12733 4215 12736
rect 4157 12727 4215 12733
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 2498 12696 2504 12708
rect 1964 12668 2504 12696
rect 1964 12640 1992 12668
rect 2498 12656 2504 12668
rect 2556 12656 2562 12708
rect 3605 12699 3663 12705
rect 3605 12665 3617 12699
rect 3651 12665 3663 12699
rect 4540 12696 4568 12724
rect 5350 12696 5356 12708
rect 4540 12668 5356 12696
rect 3605 12659 3663 12665
rect 1946 12588 1952 12640
rect 2004 12588 2010 12640
rect 2130 12588 2136 12640
rect 2188 12628 2194 12640
rect 3620 12628 3648 12659
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 5534 12656 5540 12708
rect 5592 12696 5598 12708
rect 5994 12696 6000 12708
rect 5592 12668 6000 12696
rect 5592 12656 5598 12668
rect 5994 12656 6000 12668
rect 6052 12656 6058 12708
rect 4522 12628 4528 12640
rect 2188 12600 4528 12628
rect 2188 12588 2194 12600
rect 4522 12588 4528 12600
rect 4580 12588 4586 12640
rect 5813 12631 5871 12637
rect 5813 12597 5825 12631
rect 5859 12628 5871 12631
rect 6288 12628 6316 12872
rect 7558 12860 7564 12872
rect 7616 12860 7622 12912
rect 8478 12860 8484 12912
rect 8536 12900 8542 12912
rect 9766 12900 9772 12912
rect 8536 12872 9772 12900
rect 8536 12860 8542 12872
rect 9766 12860 9772 12872
rect 9824 12860 9830 12912
rect 9858 12860 9864 12912
rect 9916 12900 9922 12912
rect 11624 12900 11652 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 12250 12968 12256 12980
rect 11977 12931 12035 12937
rect 12084 12940 12256 12968
rect 9916 12872 11652 12900
rect 11885 12903 11943 12909
rect 9916 12860 9922 12872
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 12084 12900 12112 12940
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 12713 12971 12771 12977
rect 12713 12937 12725 12971
rect 12759 12937 12771 12971
rect 12713 12931 12771 12937
rect 11931 12872 12112 12900
rect 12728 12900 12756 12931
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 13081 12971 13139 12977
rect 13081 12968 13093 12971
rect 12860 12940 13093 12968
rect 12860 12928 12866 12940
rect 13081 12937 13093 12940
rect 13127 12937 13139 12971
rect 15194 12968 15200 12980
rect 13081 12931 13139 12937
rect 13786 12940 15200 12968
rect 12728 12872 12940 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12832 6423 12835
rect 7742 12832 7748 12844
rect 6411 12804 7748 12832
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 7834 12792 7840 12844
rect 7892 12832 7898 12844
rect 7892 12804 7937 12832
rect 7892 12792 7898 12804
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 8904 12804 9413 12832
rect 8904 12792 8910 12804
rect 9401 12801 9413 12804
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 9950 12792 9956 12844
rect 10008 12838 10014 12844
rect 10137 12838 10195 12841
rect 10008 12835 10195 12838
rect 10008 12810 10149 12835
rect 10008 12792 10014 12810
rect 10137 12801 10149 12810
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 10318 12792 10324 12844
rect 10376 12832 10382 12844
rect 10594 12832 10600 12844
rect 10376 12804 10600 12832
rect 10376 12792 10382 12804
rect 10594 12792 10600 12804
rect 10652 12792 10658 12844
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10744 12804 10793 12832
rect 10744 12792 10750 12804
rect 10781 12801 10793 12804
rect 10827 12801 10839 12835
rect 10962 12832 10968 12844
rect 10923 12804 10968 12832
rect 10781 12795 10839 12801
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 11388 12804 12204 12832
rect 11388 12792 11394 12804
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 7098 12764 7104 12776
rect 6687 12736 7104 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 7098 12724 7104 12736
rect 7156 12764 7162 12776
rect 7466 12764 7472 12776
rect 7156 12736 7472 12764
rect 7156 12724 7162 12736
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 9214 12764 9220 12776
rect 7760 12736 9220 12764
rect 6362 12656 6368 12708
rect 6420 12696 6426 12708
rect 7760 12696 7788 12736
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 9490 12724 9496 12776
rect 9548 12764 9554 12776
rect 9548 12736 10824 12764
rect 9548 12724 9554 12736
rect 6420 12668 7788 12696
rect 6420 12656 6426 12668
rect 7834 12656 7840 12708
rect 7892 12696 7898 12708
rect 7892 12668 8984 12696
rect 7892 12656 7898 12668
rect 5859 12600 6316 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 8846 12628 8852 12640
rect 6604 12600 8852 12628
rect 6604 12588 6610 12600
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 8956 12628 8984 12668
rect 9306 12656 9312 12708
rect 9364 12696 9370 12708
rect 10796 12705 10824 12736
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 12069 12767 12127 12773
rect 12069 12764 12081 12767
rect 10928 12736 12081 12764
rect 10928 12724 10934 12736
rect 12069 12733 12081 12736
rect 12115 12733 12127 12767
rect 12176 12764 12204 12804
rect 12526 12792 12532 12844
rect 12584 12832 12590 12844
rect 12802 12832 12808 12844
rect 12584 12804 12808 12832
rect 12584 12792 12590 12804
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 12912 12832 12940 12872
rect 12986 12860 12992 12912
rect 13044 12900 13050 12912
rect 13446 12900 13452 12912
rect 13044 12872 13452 12900
rect 13044 12860 13050 12872
rect 13446 12860 13452 12872
rect 13504 12860 13510 12912
rect 13786 12832 13814 12940
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 15470 12968 15476 12980
rect 15431 12940 15476 12968
rect 15470 12928 15476 12940
rect 15528 12968 15534 12980
rect 15654 12968 15660 12980
rect 15528 12940 15660 12968
rect 15528 12928 15534 12940
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 13998 12860 14004 12912
rect 14056 12900 14062 12912
rect 14277 12903 14335 12909
rect 14277 12900 14289 12903
rect 14056 12872 14289 12900
rect 14056 12860 14062 12872
rect 14277 12869 14289 12872
rect 14323 12869 14335 12903
rect 14277 12863 14335 12869
rect 12912 12804 13814 12832
rect 14090 12792 14096 12844
rect 14148 12832 14154 12844
rect 14369 12835 14427 12841
rect 14148 12804 14193 12832
rect 14148 12792 14154 12804
rect 14369 12801 14381 12835
rect 14415 12832 14427 12835
rect 14642 12832 14648 12844
rect 14415 12804 14648 12832
rect 14415 12801 14427 12804
rect 14369 12795 14427 12801
rect 14642 12792 14648 12804
rect 14700 12792 14706 12844
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 15289 12835 15347 12841
rect 15289 12832 15301 12835
rect 14884 12804 15301 12832
rect 14884 12792 14890 12804
rect 15289 12801 15301 12804
rect 15335 12801 15347 12835
rect 15289 12795 15347 12801
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 15565 12835 15623 12841
rect 15565 12832 15577 12835
rect 15436 12804 15577 12832
rect 15436 12792 15442 12804
rect 15565 12801 15577 12804
rect 15611 12801 15623 12835
rect 15565 12795 15623 12801
rect 13173 12767 13231 12773
rect 13173 12764 13185 12767
rect 12176 12736 13185 12764
rect 12069 12727 12127 12733
rect 13173 12733 13185 12736
rect 13219 12733 13231 12767
rect 13173 12727 13231 12733
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 16298 12764 16304 12776
rect 13311 12736 16304 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 10781 12699 10839 12705
rect 9364 12668 10456 12696
rect 9364 12656 9370 12668
rect 9490 12628 9496 12640
rect 8956 12600 9496 12628
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 10229 12631 10287 12637
rect 10229 12597 10241 12631
rect 10275 12628 10287 12631
rect 10318 12628 10324 12640
rect 10275 12600 10324 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 10428 12628 10456 12668
rect 10781 12665 10793 12699
rect 10827 12665 10839 12699
rect 10781 12659 10839 12665
rect 11790 12656 11796 12708
rect 11848 12696 11854 12708
rect 12526 12696 12532 12708
rect 11848 12668 12532 12696
rect 11848 12656 11854 12668
rect 12526 12656 12532 12668
rect 12584 12696 12590 12708
rect 12986 12696 12992 12708
rect 12584 12668 12992 12696
rect 12584 12656 12590 12668
rect 12986 12656 12992 12668
rect 13044 12656 13050 12708
rect 12434 12628 12440 12640
rect 10428 12600 12440 12628
rect 12434 12588 12440 12600
rect 12492 12628 12498 12640
rect 13280 12628 13308 12727
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 13998 12656 14004 12708
rect 14056 12696 14062 12708
rect 14056 12668 14872 12696
rect 14056 12656 14062 12668
rect 12492 12600 13308 12628
rect 12492 12588 12498 12600
rect 13354 12588 13360 12640
rect 13412 12628 13418 12640
rect 13814 12628 13820 12640
rect 13412 12600 13820 12628
rect 13412 12588 13418 12600
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 13909 12631 13967 12637
rect 13909 12597 13921 12631
rect 13955 12628 13967 12631
rect 14090 12628 14096 12640
rect 13955 12600 14096 12628
rect 13955 12597 13967 12600
rect 13909 12591 13967 12597
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 14458 12588 14464 12640
rect 14516 12628 14522 12640
rect 14734 12628 14740 12640
rect 14516 12600 14740 12628
rect 14516 12588 14522 12600
rect 14734 12588 14740 12600
rect 14792 12588 14798 12640
rect 14844 12628 14872 12668
rect 15105 12631 15163 12637
rect 15105 12628 15117 12631
rect 14844 12600 15117 12628
rect 15105 12597 15117 12600
rect 15151 12597 15163 12631
rect 15105 12591 15163 12597
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 15746 12628 15752 12640
rect 15252 12600 15752 12628
rect 15252 12588 15258 12600
rect 15746 12588 15752 12600
rect 15804 12588 15810 12640
rect 1104 12538 16836 12560
rect 1104 12486 2924 12538
rect 2976 12486 2988 12538
rect 3040 12486 3052 12538
rect 3104 12486 3116 12538
rect 3168 12486 3180 12538
rect 3232 12486 6872 12538
rect 6924 12486 6936 12538
rect 6988 12486 7000 12538
rect 7052 12486 7064 12538
rect 7116 12486 7128 12538
rect 7180 12486 10820 12538
rect 10872 12486 10884 12538
rect 10936 12486 10948 12538
rect 11000 12486 11012 12538
rect 11064 12486 11076 12538
rect 11128 12486 14768 12538
rect 14820 12486 14832 12538
rect 14884 12486 14896 12538
rect 14948 12486 14960 12538
rect 15012 12486 15024 12538
rect 15076 12486 16836 12538
rect 1104 12464 16836 12486
rect 2038 12384 2044 12436
rect 2096 12424 2102 12436
rect 4154 12424 4160 12436
rect 2096 12396 4160 12424
rect 2096 12384 2102 12396
rect 4154 12384 4160 12396
rect 4212 12424 4218 12436
rect 5629 12427 5687 12433
rect 4212 12396 4384 12424
rect 4212 12384 4218 12396
rect 290 12316 296 12368
rect 348 12356 354 12368
rect 348 12328 1624 12356
rect 348 12316 354 12328
rect 934 12248 940 12300
rect 992 12288 998 12300
rect 1596 12297 1624 12328
rect 3050 12316 3056 12368
rect 3108 12356 3114 12368
rect 3418 12356 3424 12368
rect 3108 12328 3424 12356
rect 3108 12316 3114 12328
rect 3418 12316 3424 12328
rect 3476 12316 3482 12368
rect 3602 12316 3608 12368
rect 3660 12356 3666 12368
rect 4356 12356 4384 12396
rect 5629 12393 5641 12427
rect 5675 12424 5687 12427
rect 8662 12424 8668 12436
rect 5675 12396 8668 12424
rect 5675 12393 5687 12396
rect 5629 12387 5687 12393
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 9033 12427 9091 12433
rect 9033 12393 9045 12427
rect 9079 12424 9091 12427
rect 9306 12424 9312 12436
rect 9079 12396 9312 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 9306 12384 9312 12396
rect 9364 12424 9370 12436
rect 11330 12424 11336 12436
rect 9364 12396 11336 12424
rect 9364 12384 9370 12396
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 11440 12396 12940 12424
rect 3660 12328 4088 12356
rect 4356 12328 4568 12356
rect 3660 12316 3666 12328
rect 1397 12291 1455 12297
rect 1397 12288 1409 12291
rect 992 12260 1409 12288
rect 992 12248 998 12260
rect 1397 12257 1409 12260
rect 1443 12257 1455 12291
rect 1397 12251 1455 12257
rect 1581 12291 1639 12297
rect 1581 12257 1593 12291
rect 1627 12257 1639 12291
rect 1581 12251 1639 12257
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12288 2099 12291
rect 2130 12288 2136 12300
rect 2087 12260 2136 12288
rect 2087 12257 2099 12260
rect 2041 12251 2099 12257
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 2455 12291 2513 12297
rect 2455 12257 2467 12291
rect 2501 12288 2513 12291
rect 3142 12288 3148 12300
rect 2501 12260 3148 12288
rect 2501 12257 2513 12260
rect 2455 12251 2513 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 3878 12248 3884 12300
rect 3936 12288 3942 12300
rect 3973 12291 4031 12297
rect 3973 12288 3985 12291
rect 3936 12260 3985 12288
rect 3936 12248 3942 12260
rect 3973 12257 3985 12260
rect 4019 12257 4031 12291
rect 4060 12288 4088 12328
rect 4430 12288 4436 12300
rect 4060 12260 4436 12288
rect 3973 12251 4031 12257
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 4540 12288 4568 12328
rect 7006 12316 7012 12368
rect 7064 12356 7070 12368
rect 9674 12356 9680 12368
rect 7064 12328 9680 12356
rect 7064 12316 7070 12328
rect 9674 12316 9680 12328
rect 9732 12316 9738 12368
rect 11440 12356 11468 12396
rect 12912 12365 12940 12396
rect 13170 12384 13176 12436
rect 13228 12424 13234 12436
rect 13998 12424 14004 12436
rect 13228 12396 14004 12424
rect 13228 12384 13234 12396
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14148 12396 15056 12424
rect 14148 12384 14154 12396
rect 10888 12328 11468 12356
rect 12897 12359 12955 12365
rect 10888 12300 10916 12328
rect 12897 12325 12909 12359
rect 12943 12325 12955 12359
rect 12897 12319 12955 12325
rect 4709 12291 4767 12297
rect 4709 12288 4721 12291
rect 4540 12260 4721 12288
rect 4709 12257 4721 12260
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 4982 12248 4988 12300
rect 5040 12288 5046 12300
rect 5040 12260 5580 12288
rect 5040 12248 5046 12260
rect 2314 12180 2320 12232
rect 2372 12220 2378 12232
rect 2590 12220 2596 12232
rect 2372 12192 2417 12220
rect 2551 12192 2596 12220
rect 2372 12180 2378 12192
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 3789 12223 3847 12229
rect 3789 12220 3801 12223
rect 3476 12192 3801 12220
rect 3476 12180 3482 12192
rect 3789 12189 3801 12192
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 4798 12180 4804 12232
rect 4856 12229 4862 12232
rect 4856 12223 4884 12229
rect 4872 12189 4884 12223
rect 4856 12183 4884 12189
rect 4856 12180 4862 12183
rect 3237 12155 3295 12161
rect 3237 12121 3249 12155
rect 3283 12152 3295 12155
rect 3878 12152 3884 12164
rect 3283 12124 3884 12152
rect 3283 12121 3295 12124
rect 3237 12115 3295 12121
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 5552 12152 5580 12260
rect 6730 12248 6736 12300
rect 6788 12288 6794 12300
rect 6788 12260 9820 12288
rect 6788 12248 6794 12260
rect 6914 12220 6920 12232
rect 6564 12192 6920 12220
rect 6564 12152 6592 12192
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 8018 12180 8024 12232
rect 8076 12220 8082 12232
rect 9217 12223 9275 12229
rect 9217 12220 9229 12223
rect 8076 12192 9229 12220
rect 8076 12180 8082 12192
rect 9217 12189 9229 12192
rect 9263 12189 9275 12223
rect 9674 12220 9680 12232
rect 9635 12192 9680 12220
rect 9217 12183 9275 12189
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 9792 12220 9820 12260
rect 10870 12248 10876 12300
rect 10928 12248 10934 12300
rect 12912 12288 12940 12319
rect 13078 12316 13084 12368
rect 13136 12356 13142 12368
rect 13357 12359 13415 12365
rect 13357 12356 13369 12359
rect 13136 12328 13369 12356
rect 13136 12316 13142 12328
rect 13357 12325 13369 12328
rect 13403 12325 13415 12359
rect 13357 12319 13415 12325
rect 13446 12316 13452 12368
rect 13504 12356 13510 12368
rect 14642 12356 14648 12368
rect 13504 12328 14648 12356
rect 13504 12316 13510 12328
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 15028 12356 15056 12396
rect 15102 12384 15108 12436
rect 15160 12424 15166 12436
rect 15378 12424 15384 12436
rect 15160 12396 15384 12424
rect 15160 12384 15166 12396
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 15654 12356 15660 12368
rect 15028 12328 15660 12356
rect 15654 12316 15660 12328
rect 15712 12316 15718 12368
rect 11440 12260 11652 12288
rect 12912 12260 13768 12288
rect 11440 12220 11468 12260
rect 9792 12192 11468 12220
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12189 11575 12223
rect 11624 12220 11652 12260
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 11624 12192 13553 12220
rect 11517 12183 11575 12189
rect 13541 12189 13553 12192
rect 13587 12220 13599 12223
rect 13630 12220 13636 12232
rect 13587 12192 13636 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 5552 12124 6592 12152
rect 6641 12155 6699 12161
rect 6641 12121 6653 12155
rect 6687 12152 6699 12155
rect 7006 12152 7012 12164
rect 6687 12124 7012 12152
rect 6687 12121 6699 12124
rect 6641 12115 6699 12121
rect 7006 12112 7012 12124
rect 7064 12112 7070 12164
rect 8110 12112 8116 12164
rect 8168 12152 8174 12164
rect 9950 12161 9956 12164
rect 8168 12124 8984 12152
rect 8168 12112 8174 12124
rect 2682 12044 2688 12096
rect 2740 12084 2746 12096
rect 5902 12084 5908 12096
rect 2740 12056 5908 12084
rect 2740 12044 2746 12056
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 6270 12044 6276 12096
rect 6328 12084 6334 12096
rect 6822 12084 6828 12096
rect 6328 12056 6828 12084
rect 6328 12044 6334 12056
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 7929 12087 7987 12093
rect 7929 12084 7941 12087
rect 7248 12056 7941 12084
rect 7248 12044 7254 12056
rect 7929 12053 7941 12056
rect 7975 12053 7987 12087
rect 7929 12047 7987 12053
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8478 12084 8484 12096
rect 8260 12056 8484 12084
rect 8260 12044 8266 12056
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 8956 12084 8984 12124
rect 9944 12115 9956 12161
rect 10008 12152 10014 12164
rect 11532 12152 11560 12183
rect 13630 12180 13636 12192
rect 13688 12180 13694 12232
rect 13740 12220 13768 12260
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 14090 12288 14096 12300
rect 13964 12260 14096 12288
rect 13964 12248 13970 12260
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 14366 12288 14372 12300
rect 14279 12260 14372 12288
rect 14292 12229 14320 12260
rect 14366 12248 14372 12260
rect 14424 12288 14430 12300
rect 14424 12260 15148 12288
rect 14424 12248 14430 12260
rect 15120 12232 15148 12260
rect 14277 12223 14335 12229
rect 13740 12192 14228 12220
rect 10008 12124 10044 12152
rect 10144 12124 11560 12152
rect 11784 12155 11842 12161
rect 9950 12112 9956 12115
rect 10008 12112 10014 12124
rect 10144 12084 10172 12124
rect 11784 12121 11796 12155
rect 11830 12152 11842 12155
rect 14093 12155 14151 12161
rect 14093 12152 14105 12155
rect 11830 12124 14105 12152
rect 11830 12121 11842 12124
rect 11784 12115 11842 12121
rect 14093 12121 14105 12124
rect 14139 12121 14151 12155
rect 14200 12152 14228 12192
rect 14277 12189 14289 12223
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12220 14611 12223
rect 14642 12220 14648 12232
rect 14599 12192 14648 12220
rect 14599 12189 14611 12192
rect 14553 12183 14611 12189
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 15102 12180 15108 12232
rect 15160 12220 15166 12232
rect 15197 12223 15255 12229
rect 15197 12220 15209 12223
rect 15160 12192 15209 12220
rect 15160 12180 15166 12192
rect 15197 12189 15209 12192
rect 15243 12189 15255 12223
rect 15197 12183 15255 12189
rect 15470 12180 15476 12232
rect 15528 12220 15534 12232
rect 15930 12220 15936 12232
rect 15528 12192 15573 12220
rect 15891 12192 15936 12220
rect 15528 12180 15534 12192
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 14461 12155 14519 12161
rect 14461 12152 14473 12155
rect 14200 12124 14473 12152
rect 14093 12115 14151 12121
rect 14461 12121 14473 12124
rect 14507 12121 14519 12155
rect 14461 12115 14519 12121
rect 14918 12112 14924 12164
rect 14976 12152 14982 12164
rect 14976 12124 15424 12152
rect 14976 12112 14982 12124
rect 11054 12084 11060 12096
rect 8956 12056 10172 12084
rect 11015 12056 11060 12084
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 12894 12084 12900 12096
rect 11204 12056 12900 12084
rect 11204 12044 11210 12056
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 15396 12093 15424 12124
rect 15562 12112 15568 12164
rect 15620 12152 15626 12164
rect 15620 12124 15792 12152
rect 15620 12112 15626 12124
rect 15013 12087 15071 12093
rect 15013 12084 15025 12087
rect 13320 12056 15025 12084
rect 13320 12044 13326 12056
rect 15013 12053 15025 12056
rect 15059 12053 15071 12087
rect 15013 12047 15071 12053
rect 15381 12087 15439 12093
rect 15381 12053 15393 12087
rect 15427 12053 15439 12087
rect 15764 12084 15792 12124
rect 15930 12084 15936 12096
rect 15764 12056 15936 12084
rect 15381 12047 15439 12053
rect 15930 12044 15936 12056
rect 15988 12044 15994 12096
rect 16117 12087 16175 12093
rect 16117 12053 16129 12087
rect 16163 12084 16175 12087
rect 16390 12084 16396 12096
rect 16163 12056 16396 12084
rect 16163 12053 16175 12056
rect 16117 12047 16175 12053
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 1104 11994 16836 12016
rect 1104 11942 4898 11994
rect 4950 11942 4962 11994
rect 5014 11942 5026 11994
rect 5078 11942 5090 11994
rect 5142 11942 5154 11994
rect 5206 11942 8846 11994
rect 8898 11942 8910 11994
rect 8962 11942 8974 11994
rect 9026 11942 9038 11994
rect 9090 11942 9102 11994
rect 9154 11942 12794 11994
rect 12846 11942 12858 11994
rect 12910 11942 12922 11994
rect 12974 11942 12986 11994
rect 13038 11942 13050 11994
rect 13102 11942 16836 11994
rect 1104 11920 16836 11942
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 2958 11880 2964 11892
rect 2832 11852 2964 11880
rect 2832 11840 2838 11852
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 3418 11840 3424 11892
rect 3476 11880 3482 11892
rect 4706 11880 4712 11892
rect 3476 11852 4568 11880
rect 4667 11852 4712 11880
rect 3476 11840 3482 11852
rect 4540 11812 4568 11852
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5132 11852 5672 11880
rect 5132 11840 5138 11852
rect 4540 11784 5488 11812
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11744 1642 11756
rect 2130 11744 2136 11756
rect 1636 11716 2136 11744
rect 1636 11704 1642 11716
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11744 3111 11747
rect 3234 11744 3240 11756
rect 3099 11716 3240 11744
rect 3099 11713 3111 11716
rect 3053 11707 3111 11713
rect 3234 11704 3240 11716
rect 3292 11704 3298 11756
rect 4062 11744 4068 11756
rect 4023 11716 4068 11744
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 5166 11744 5172 11756
rect 5127 11716 5172 11744
rect 5166 11704 5172 11716
rect 5224 11704 5230 11756
rect 5460 11753 5488 11784
rect 5644 11753 5672 11852
rect 6472 11852 8340 11880
rect 6472 11756 6500 11852
rect 8110 11812 8116 11824
rect 6564 11784 8116 11812
rect 5445 11747 5503 11753
rect 5445 11713 5457 11747
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 1857 11679 1915 11685
rect 1857 11645 1869 11679
rect 1903 11676 1915 11679
rect 2222 11676 2228 11688
rect 1903 11648 2228 11676
rect 1903 11645 1915 11648
rect 1857 11639 1915 11645
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 2869 11679 2927 11685
rect 2869 11645 2881 11679
rect 2915 11645 2927 11679
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 2869 11639 2927 11645
rect 3620 11648 3801 11676
rect 2884 11608 2912 11639
rect 3050 11608 3056 11620
rect 2884 11580 3056 11608
rect 3050 11568 3056 11580
rect 3108 11568 3114 11620
rect 3510 11608 3516 11620
rect 3471 11580 3516 11608
rect 3510 11568 3516 11580
rect 3568 11568 3574 11620
rect 382 11500 388 11552
rect 440 11540 446 11552
rect 2038 11540 2044 11552
rect 440 11512 2044 11540
rect 440 11500 446 11512
rect 2038 11500 2044 11512
rect 2096 11500 2102 11552
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 3620 11540 3648 11648
rect 3789 11645 3801 11648
rect 3835 11645 3847 11679
rect 3789 11639 3847 11645
rect 3927 11679 3985 11685
rect 3927 11645 3939 11679
rect 3973 11676 3985 11679
rect 3973 11648 5396 11676
rect 3973 11645 3985 11648
rect 3927 11639 3985 11645
rect 5166 11540 5172 11552
rect 2372 11512 5172 11540
rect 2372 11500 2378 11512
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 5368 11540 5396 11648
rect 5460 11608 5488 11707
rect 5718 11704 5724 11756
rect 5776 11744 5782 11756
rect 6454 11744 6460 11756
rect 5776 11716 6460 11744
rect 5776 11704 5782 11716
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 6564 11753 6592 11784
rect 8110 11772 8116 11784
rect 8168 11772 8174 11824
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 6816 11747 6874 11753
rect 6816 11713 6828 11747
rect 6862 11744 6874 11747
rect 8202 11744 8208 11756
rect 6862 11716 8208 11744
rect 6862 11713 6874 11716
rect 6816 11707 6874 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 8312 11744 8340 11852
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 9677 11883 9735 11889
rect 9677 11880 9689 11883
rect 9640 11852 9689 11880
rect 9640 11840 9646 11852
rect 9677 11849 9689 11852
rect 9723 11849 9735 11883
rect 9677 11843 9735 11849
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 10502 11880 10508 11892
rect 10376 11852 10508 11880
rect 10376 11840 10382 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 10652 11852 10697 11880
rect 10652 11840 10658 11852
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 11330 11880 11336 11892
rect 10836 11852 11336 11880
rect 10836 11840 10842 11852
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 11422 11840 11428 11892
rect 11480 11880 11486 11892
rect 13262 11880 13268 11892
rect 11480 11852 13268 11880
rect 11480 11840 11486 11852
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13722 11840 13728 11892
rect 13780 11840 13786 11892
rect 13909 11883 13967 11889
rect 13909 11849 13921 11883
rect 13955 11849 13967 11883
rect 13909 11843 13967 11849
rect 8389 11815 8447 11821
rect 8389 11781 8401 11815
rect 8435 11812 8447 11815
rect 13170 11812 13176 11824
rect 8435 11784 13176 11812
rect 8435 11781 8447 11784
rect 8389 11775 8447 11781
rect 13170 11772 13176 11784
rect 13228 11772 13234 11824
rect 13446 11772 13452 11824
rect 13504 11772 13510 11824
rect 8312 11716 9076 11744
rect 5810 11676 5816 11688
rect 5771 11648 5816 11676
rect 5810 11636 5816 11648
rect 5868 11636 5874 11688
rect 9048 11676 9076 11716
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 9180 11716 10793 11744
rect 9180 11704 9186 11716
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11773 11747 11831 11753
rect 11773 11744 11785 11747
rect 11664 11716 11785 11744
rect 11664 11704 11670 11716
rect 11773 11713 11785 11716
rect 11819 11713 11831 11747
rect 11773 11707 11831 11713
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12124 11716 12572 11744
rect 12124 11704 12130 11716
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 9048 11648 11529 11676
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 6270 11608 6276 11620
rect 5460 11580 6276 11608
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 8386 11568 8392 11620
rect 8444 11608 8450 11620
rect 12544 11608 12572 11716
rect 12710 11704 12716 11756
rect 12768 11744 12774 11756
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 12768 11716 13369 11744
rect 12768 11704 12774 11716
rect 13357 11713 13369 11716
rect 13403 11713 13415 11747
rect 13357 11707 13415 11713
rect 13464 11744 13492 11772
rect 13740 11753 13768 11840
rect 13924 11812 13952 11843
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 15381 11883 15439 11889
rect 15381 11880 15393 11883
rect 15344 11852 15393 11880
rect 15344 11840 15350 11852
rect 15381 11849 15393 11852
rect 15427 11849 15439 11883
rect 15381 11843 15439 11849
rect 14366 11812 14372 11824
rect 13924 11784 14372 11812
rect 14366 11772 14372 11784
rect 14424 11772 14430 11824
rect 14734 11812 14740 11824
rect 14695 11784 14740 11812
rect 14734 11772 14740 11784
rect 14792 11772 14798 11824
rect 15749 11815 15807 11821
rect 15749 11812 15761 11815
rect 14844 11784 15761 11812
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 13464 11716 13553 11744
rect 13464 11676 13492 11716
rect 13541 11713 13553 11716
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11713 13783 11747
rect 14844 11744 14872 11784
rect 15749 11781 15761 11784
rect 15795 11781 15807 11815
rect 15749 11775 15807 11781
rect 13725 11707 13783 11713
rect 14108 11716 14872 11744
rect 13188 11648 13492 11676
rect 13644 11676 13672 11707
rect 14108 11688 14136 11716
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15565 11747 15623 11753
rect 15565 11744 15577 11747
rect 15344 11716 15577 11744
rect 15344 11704 15350 11716
rect 15565 11713 15577 11716
rect 15611 11713 15623 11747
rect 15565 11707 15623 11713
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 14090 11676 14096 11688
rect 13644 11648 14096 11676
rect 12897 11611 12955 11617
rect 12897 11608 12909 11611
rect 8444 11580 11560 11608
rect 12544 11580 12909 11608
rect 8444 11568 8450 11580
rect 5626 11540 5632 11552
rect 5368 11512 5632 11540
rect 5626 11500 5632 11512
rect 5684 11540 5690 11552
rect 7466 11540 7472 11552
rect 5684 11512 7472 11540
rect 5684 11500 5690 11512
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 7929 11543 7987 11549
rect 7929 11509 7941 11543
rect 7975 11540 7987 11543
rect 10226 11540 10232 11552
rect 7975 11512 10232 11540
rect 7975 11509 7987 11512
rect 7929 11503 7987 11509
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 11532 11540 11560 11580
rect 12897 11577 12909 11580
rect 12943 11577 12955 11611
rect 12897 11571 12955 11577
rect 13188 11540 13216 11648
rect 14090 11636 14096 11648
rect 14148 11636 14154 11688
rect 14642 11636 14648 11688
rect 14700 11676 14706 11688
rect 15856 11676 15884 11707
rect 14700 11648 15884 11676
rect 14700 11636 14706 11648
rect 13262 11568 13268 11620
rect 13320 11608 13326 11620
rect 14369 11611 14427 11617
rect 14369 11608 14381 11611
rect 13320 11580 14381 11608
rect 13320 11568 13326 11580
rect 14369 11577 14381 11580
rect 14415 11577 14427 11611
rect 14369 11571 14427 11577
rect 14921 11611 14979 11617
rect 14921 11577 14933 11611
rect 14967 11608 14979 11611
rect 14967 11580 16896 11608
rect 14967 11577 14979 11580
rect 14921 11571 14979 11577
rect 11532 11512 13216 11540
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14182 11540 14188 11552
rect 13872 11512 14188 11540
rect 13872 11500 13878 11512
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 14759 11543 14817 11549
rect 14759 11509 14771 11543
rect 14805 11540 14817 11543
rect 16114 11540 16120 11552
rect 14805 11512 16120 11540
rect 14805 11509 14817 11512
rect 14759 11503 14817 11509
rect 16114 11500 16120 11512
rect 16172 11500 16178 11552
rect 1104 11450 16836 11472
rect 1104 11398 2924 11450
rect 2976 11398 2988 11450
rect 3040 11398 3052 11450
rect 3104 11398 3116 11450
rect 3168 11398 3180 11450
rect 3232 11398 6872 11450
rect 6924 11398 6936 11450
rect 6988 11398 7000 11450
rect 7052 11398 7064 11450
rect 7116 11398 7128 11450
rect 7180 11398 10820 11450
rect 10872 11398 10884 11450
rect 10936 11398 10948 11450
rect 11000 11398 11012 11450
rect 11064 11398 11076 11450
rect 11128 11398 14768 11450
rect 14820 11398 14832 11450
rect 14884 11398 14896 11450
rect 14948 11398 14960 11450
rect 15012 11398 15024 11450
rect 15076 11398 16836 11450
rect 1104 11376 16836 11398
rect 16868 11404 16896 11580
rect 16868 11376 16988 11404
rect 10778 11336 10784 11348
rect 3160 11308 10784 11336
rect 1489 11203 1547 11209
rect 1489 11169 1501 11203
rect 1535 11200 1547 11203
rect 2958 11200 2964 11212
rect 1535 11172 2964 11200
rect 1535 11169 1547 11172
rect 1489 11163 1547 11169
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 3160 11132 3188 11308
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 11974 11336 11980 11348
rect 11808 11308 11980 11336
rect 3237 11271 3295 11277
rect 3237 11237 3249 11271
rect 3283 11268 3295 11271
rect 4062 11268 4068 11280
rect 3283 11240 4068 11268
rect 3283 11237 3295 11240
rect 3237 11231 3295 11237
rect 4062 11228 4068 11240
rect 4120 11228 4126 11280
rect 4172 11240 4568 11268
rect 4172 11200 4200 11240
rect 3804 11172 4200 11200
rect 3804 11141 3832 11172
rect 4246 11160 4252 11212
rect 4304 11200 4310 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4304 11172 4445 11200
rect 4304 11160 4310 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4540 11200 4568 11240
rect 5902 11228 5908 11280
rect 5960 11268 5966 11280
rect 6181 11271 6239 11277
rect 6181 11268 6193 11271
rect 5960 11240 6193 11268
rect 5960 11228 5966 11240
rect 6181 11237 6193 11240
rect 6227 11237 6239 11271
rect 6181 11231 6239 11237
rect 6270 11228 6276 11280
rect 6328 11268 6334 11280
rect 6454 11268 6460 11280
rect 6328 11240 6460 11268
rect 6328 11228 6334 11240
rect 6454 11228 6460 11240
rect 6512 11228 6518 11280
rect 7466 11268 7472 11280
rect 7300 11240 7472 11268
rect 7300 11200 7328 11240
rect 7466 11228 7472 11240
rect 7524 11228 7530 11280
rect 10134 11228 10140 11280
rect 10192 11268 10198 11280
rect 10318 11268 10324 11280
rect 10192 11240 10324 11268
rect 10192 11228 10198 11240
rect 10318 11228 10324 11240
rect 10376 11228 10382 11280
rect 10410 11228 10416 11280
rect 10468 11268 10474 11280
rect 10594 11268 10600 11280
rect 10468 11240 10600 11268
rect 10468 11228 10474 11240
rect 10594 11228 10600 11240
rect 10652 11228 10658 11280
rect 4540 11172 7328 11200
rect 4433 11163 4491 11169
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 7834 11200 7840 11212
rect 7432 11172 7840 11200
rect 7432 11160 7438 11172
rect 7834 11160 7840 11172
rect 7892 11160 7898 11212
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8720 11172 8953 11200
rect 8720 11160 8726 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 2898 11104 3188 11132
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 8389 11135 8447 11141
rect 7156 11104 8340 11132
rect 7156 11092 7162 11104
rect 1765 11067 1823 11073
rect 1765 11033 1777 11067
rect 1811 11064 1823 11067
rect 1854 11064 1860 11076
rect 1811 11036 1860 11064
rect 1811 11033 1823 11036
rect 1765 11027 1823 11033
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 3418 11024 3424 11076
rect 3476 11064 3482 11076
rect 3881 11067 3939 11073
rect 3881 11064 3893 11067
rect 3476 11036 3893 11064
rect 3476 11024 3482 11036
rect 3881 11033 3893 11036
rect 3927 11033 3939 11067
rect 3881 11027 3939 11033
rect 4154 11024 4160 11076
rect 4212 11064 4218 11076
rect 4709 11067 4767 11073
rect 4709 11064 4721 11067
rect 4212 11036 4721 11064
rect 4212 11024 4218 11036
rect 4709 11033 4721 11036
rect 4755 11033 4767 11067
rect 6454 11064 6460 11076
rect 5934 11036 6460 11064
rect 4709 11027 4767 11033
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 6641 11067 6699 11073
rect 6641 11033 6653 11067
rect 6687 11064 6699 11067
rect 7834 11064 7840 11076
rect 6687 11036 7840 11064
rect 6687 11033 6699 11036
rect 6641 11027 6699 11033
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 8312 11064 8340 11104
rect 8389 11101 8401 11135
rect 8435 11132 8447 11135
rect 8435 11104 9720 11132
rect 8435 11101 8447 11104
rect 8389 11095 8447 11101
rect 9692 11076 9720 11104
rect 9950 11092 9956 11144
rect 10008 11132 10014 11144
rect 10686 11132 10692 11144
rect 10008 11104 10692 11132
rect 10008 11092 10014 11104
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 11514 11132 11520 11144
rect 10827 11104 11520 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 9030 11064 9036 11076
rect 8312 11036 9036 11064
rect 9030 11024 9036 11036
rect 9088 11024 9094 11076
rect 9208 11067 9266 11073
rect 9208 11033 9220 11067
rect 9254 11064 9266 11067
rect 9582 11064 9588 11076
rect 9254 11036 9588 11064
rect 9254 11033 9266 11036
rect 9208 11027 9266 11033
rect 9582 11024 9588 11036
rect 9640 11024 9646 11076
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 10870 11064 10876 11076
rect 9732 11036 10876 11064
rect 9732 11024 9738 11036
rect 10870 11024 10876 11036
rect 10928 11024 10934 11076
rect 11048 11067 11106 11073
rect 11048 11033 11060 11067
rect 11094 11064 11106 11067
rect 11238 11064 11244 11076
rect 11094 11036 11244 11064
rect 11094 11033 11106 11036
rect 11048 11027 11106 11033
rect 11238 11024 11244 11036
rect 11296 11024 11302 11076
rect 11422 11024 11428 11076
rect 11480 11064 11486 11076
rect 11808 11064 11836 11308
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 12158 11296 12164 11348
rect 12216 11336 12222 11348
rect 12216 11308 12261 11336
rect 12216 11296 12222 11308
rect 12618 11296 12624 11348
rect 12676 11336 12682 11348
rect 12802 11336 12808 11348
rect 12676 11308 12808 11336
rect 12676 11296 12682 11308
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 13004 11308 13553 11336
rect 13004 11200 13032 11308
rect 13541 11305 13553 11308
rect 13587 11305 13599 11339
rect 13541 11299 13599 11305
rect 13628 11308 13952 11336
rect 13170 11228 13176 11280
rect 13228 11268 13234 11280
rect 13628 11268 13656 11308
rect 13228 11240 13656 11268
rect 13924 11268 13952 11308
rect 14090 11296 14096 11348
rect 14148 11336 14154 11348
rect 15194 11336 15200 11348
rect 14148 11308 15200 11336
rect 14148 11296 14154 11308
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 16114 11296 16120 11348
rect 16172 11336 16178 11348
rect 16850 11336 16856 11348
rect 16172 11308 16856 11336
rect 16172 11296 16178 11308
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 14645 11271 14703 11277
rect 13924 11240 14412 11268
rect 13228 11228 13234 11240
rect 12268 11172 13032 11200
rect 12066 11092 12072 11144
rect 12124 11092 12130 11144
rect 12158 11092 12164 11144
rect 12216 11132 12222 11144
rect 12268 11132 12296 11172
rect 12216 11104 12296 11132
rect 12216 11092 12222 11104
rect 12802 11092 12808 11144
rect 12860 11142 12866 11144
rect 12860 11141 13032 11142
rect 12860 11135 13047 11141
rect 12860 11114 13001 11135
rect 12860 11092 12866 11114
rect 12989 11101 13001 11114
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 13078 11092 13084 11144
rect 13136 11132 13142 11144
rect 13280 11141 13308 11240
rect 13630 11160 13636 11212
rect 13688 11200 13694 11212
rect 14384 11200 14412 11240
rect 14645 11237 14657 11271
rect 14691 11268 14703 11271
rect 14918 11268 14924 11280
rect 14691 11240 14924 11268
rect 14691 11237 14703 11240
rect 14645 11231 14703 11237
rect 14918 11228 14924 11240
rect 14976 11228 14982 11280
rect 13688 11172 14320 11200
rect 14384 11172 15516 11200
rect 13688 11160 13694 11172
rect 13173 11135 13231 11141
rect 13173 11132 13185 11135
rect 13136 11104 13185 11132
rect 13136 11092 13142 11104
rect 13173 11101 13185 11104
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 13381 11135 13439 11141
rect 13381 11101 13393 11135
rect 13427 11134 13439 11135
rect 13427 11132 13552 11134
rect 13722 11132 13728 11144
rect 13427 11106 13728 11132
rect 13427 11104 13446 11106
rect 13524 11104 13728 11106
rect 13427 11101 13439 11104
rect 13381 11095 13439 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 14090 11092 14096 11144
rect 14148 11132 14154 11144
rect 14292 11141 14320 11172
rect 14277 11135 14335 11141
rect 14148 11104 14193 11132
rect 14148 11092 14154 11104
rect 14277 11101 14289 11135
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 14642 11132 14648 11144
rect 14507 11104 14648 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 15286 11132 15292 11144
rect 15247 11104 15292 11132
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 15488 11141 15516 11172
rect 16850 11160 16856 11212
rect 16908 11200 16914 11212
rect 16960 11200 16988 11376
rect 16908 11172 16988 11200
rect 16908 11160 16914 11172
rect 15473 11135 15531 11141
rect 15473 11101 15485 11135
rect 15519 11101 15531 11135
rect 15473 11095 15531 11101
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11101 15623 11135
rect 15565 11095 15623 11101
rect 11480 11036 11836 11064
rect 11480 11024 11486 11036
rect 1578 10956 1584 11008
rect 1636 10996 1642 11008
rect 2590 10996 2596 11008
rect 1636 10968 2596 10996
rect 1636 10956 1642 10968
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 3326 10956 3332 11008
rect 3384 10996 3390 11008
rect 5534 10996 5540 11008
rect 3384 10968 5540 10996
rect 3384 10956 3390 10968
rect 5534 10956 5540 10968
rect 5592 10956 5598 11008
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 9122 10996 9128 11008
rect 7340 10968 9128 10996
rect 7340 10956 7346 10968
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 9766 10956 9772 11008
rect 9824 10996 9830 11008
rect 10321 10999 10379 11005
rect 10321 10996 10333 10999
rect 9824 10968 10333 10996
rect 9824 10956 9830 10968
rect 10321 10965 10333 10968
rect 10367 10965 10379 10999
rect 10321 10959 10379 10965
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 12084 10996 12112 11092
rect 14369 11067 14427 11073
rect 14369 11064 14381 11067
rect 13740 11036 14381 11064
rect 12986 10996 12992 11008
rect 10652 10968 12992 10996
rect 10652 10956 10658 10968
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13740 10996 13768 11036
rect 14369 11033 14381 11036
rect 14415 11033 14427 11067
rect 14369 11027 14427 11033
rect 14550 11024 14556 11076
rect 14608 11064 14614 11076
rect 15580 11064 15608 11095
rect 14608 11036 15608 11064
rect 14608 11024 14614 11036
rect 13412 10968 13768 10996
rect 13412 10956 13418 10968
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 15105 10999 15163 11005
rect 15105 10996 15117 10999
rect 14240 10968 15117 10996
rect 14240 10956 14246 10968
rect 15105 10965 15117 10968
rect 15151 10965 15163 10999
rect 15105 10959 15163 10965
rect 1104 10906 16836 10928
rect 1104 10854 4898 10906
rect 4950 10854 4962 10906
rect 5014 10854 5026 10906
rect 5078 10854 5090 10906
rect 5142 10854 5154 10906
rect 5206 10854 8846 10906
rect 8898 10854 8910 10906
rect 8962 10854 8974 10906
rect 9026 10854 9038 10906
rect 9090 10854 9102 10906
rect 9154 10854 12794 10906
rect 12846 10854 12858 10906
rect 12910 10854 12922 10906
rect 12974 10854 12986 10906
rect 13038 10854 13050 10906
rect 13102 10854 16836 10906
rect 1104 10832 16836 10854
rect 1762 10792 1768 10804
rect 1723 10764 1768 10792
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 2041 10795 2099 10801
rect 2041 10761 2053 10795
rect 2087 10792 2099 10795
rect 2130 10792 2136 10804
rect 2087 10764 2136 10792
rect 2087 10761 2099 10764
rect 2041 10755 2099 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 4614 10752 4620 10804
rect 4672 10792 4678 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 4672 10764 5181 10792
rect 4672 10752 4678 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 10962 10792 10968 10804
rect 5169 10755 5227 10761
rect 7760 10764 10968 10792
rect 7760 10724 7788 10764
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 12526 10792 12532 10804
rect 11716 10764 12532 10792
rect 3910 10696 7788 10724
rect 7837 10727 7895 10733
rect 7837 10693 7849 10727
rect 7883 10724 7895 10727
rect 11716 10724 11744 10764
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 12897 10795 12955 10801
rect 12897 10761 12909 10795
rect 12943 10792 12955 10795
rect 13170 10792 13176 10804
rect 12943 10764 13176 10792
rect 12943 10761 12955 10764
rect 12897 10755 12955 10761
rect 13170 10752 13176 10764
rect 13228 10752 13234 10804
rect 14182 10792 14188 10804
rect 13464 10764 14188 10792
rect 7883 10696 11744 10724
rect 11784 10727 11842 10733
rect 7883 10693 7895 10696
rect 7837 10687 7895 10693
rect 11784 10693 11796 10727
rect 11830 10724 11842 10727
rect 13464 10724 13492 10764
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 15013 10795 15071 10801
rect 14384 10764 14944 10792
rect 11830 10696 13492 10724
rect 11830 10693 11842 10696
rect 11784 10687 11842 10693
rect 13722 10684 13728 10736
rect 13780 10724 13786 10736
rect 13780 10696 13825 10724
rect 13780 10684 13786 10696
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10656 1455 10659
rect 1762 10656 1768 10668
rect 1443 10628 1768 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 1882 10659 1940 10665
rect 1882 10625 1894 10659
rect 1928 10625 1940 10659
rect 1882 10619 1940 10625
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10656 2559 10659
rect 2547 10628 2820 10656
rect 2547 10625 2559 10628
rect 2501 10619 2559 10625
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 1673 10591 1731 10597
rect 1673 10588 1685 10591
rect 1636 10560 1685 10588
rect 1636 10548 1642 10560
rect 1673 10557 1685 10560
rect 1719 10557 1731 10591
rect 1897 10588 1925 10619
rect 2682 10588 2688 10600
rect 1897 10560 2688 10588
rect 1673 10551 1731 10557
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 2792 10588 2820 10628
rect 2866 10616 2872 10668
rect 2924 10656 2930 10668
rect 2924 10628 2969 10656
rect 2924 10616 2930 10628
rect 3694 10616 3700 10668
rect 3752 10656 3758 10668
rect 4295 10659 4353 10665
rect 4295 10656 4307 10659
rect 3752 10628 4307 10656
rect 3752 10616 3758 10628
rect 4295 10625 4307 10628
rect 4341 10625 4353 10659
rect 6641 10659 6699 10665
rect 4295 10619 4353 10625
rect 4540 10628 6596 10656
rect 4540 10588 4568 10628
rect 2792 10560 4568 10588
rect 5166 10548 5172 10600
rect 5224 10588 5230 10600
rect 5261 10591 5319 10597
rect 5261 10588 5273 10591
rect 5224 10560 5273 10588
rect 5224 10548 5230 10560
rect 5261 10557 5273 10560
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 5350 10548 5356 10600
rect 5408 10588 5414 10600
rect 6365 10591 6423 10597
rect 5408 10560 5453 10588
rect 5408 10548 5414 10560
rect 6365 10557 6377 10591
rect 6411 10557 6423 10591
rect 6568 10588 6596 10628
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 8478 10656 8484 10668
rect 6687 10628 8484 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 8478 10616 8484 10628
rect 8536 10656 8542 10668
rect 8754 10656 8760 10668
rect 8536 10628 8760 10656
rect 8536 10616 8542 10628
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10134 10656 10140 10668
rect 10008 10628 10140 10656
rect 10008 10616 10014 10628
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 11146 10656 11152 10668
rect 10244 10628 11152 10656
rect 10244 10588 10272 10628
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 12802 10616 12808 10668
rect 12860 10656 12866 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 12860 10628 13553 10656
rect 12860 10616 12866 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 13630 10616 13636 10668
rect 13688 10656 13694 10668
rect 13909 10659 13967 10665
rect 13688 10628 13732 10656
rect 13688 10616 13694 10628
rect 13909 10625 13921 10659
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 14001 10659 14059 10665
rect 14001 10625 14013 10659
rect 14047 10656 14059 10659
rect 14090 10656 14096 10668
rect 14047 10628 14096 10656
rect 14047 10625 14059 10628
rect 14001 10619 14059 10625
rect 6568 10560 10272 10588
rect 10413 10591 10471 10597
rect 6365 10551 6423 10557
rect 10413 10557 10425 10591
rect 10459 10588 10471 10591
rect 10594 10588 10600 10600
rect 10459 10560 10600 10588
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 5074 10520 5080 10532
rect 3620 10492 5080 10520
rect 934 10412 940 10464
rect 992 10452 998 10464
rect 3620 10452 3648 10492
rect 5074 10480 5080 10492
rect 5132 10480 5138 10532
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 6178 10520 6184 10532
rect 5592 10492 6184 10520
rect 5592 10480 5598 10492
rect 6178 10480 6184 10492
rect 6236 10480 6242 10532
rect 6380 10520 6408 10551
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 11514 10588 11520 10600
rect 11475 10560 11520 10588
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 13924 10588 13952 10619
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 14384 10588 14412 10764
rect 14550 10684 14556 10736
rect 14608 10724 14614 10736
rect 14645 10727 14703 10733
rect 14645 10724 14657 10727
rect 14608 10696 14657 10724
rect 14608 10684 14614 10696
rect 14645 10693 14657 10696
rect 14691 10693 14703 10727
rect 14645 10687 14703 10693
rect 14734 10684 14740 10736
rect 14792 10724 14798 10736
rect 14916 10724 14944 10764
rect 15013 10761 15025 10795
rect 15059 10792 15071 10795
rect 15286 10792 15292 10804
rect 15059 10764 15292 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 16114 10792 16120 10804
rect 15396 10764 16120 10792
rect 15396 10724 15424 10764
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 14792 10696 14837 10724
rect 14916 10696 15424 10724
rect 15841 10727 15899 10733
rect 14792 10684 14798 10696
rect 15841 10693 15853 10727
rect 15887 10724 15899 10727
rect 15887 10696 16068 10724
rect 15887 10693 15899 10696
rect 15841 10687 15899 10693
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10656 14519 10659
rect 14826 10656 14832 10668
rect 14507 10628 14688 10656
rect 14787 10628 14832 10656
rect 14507 10625 14519 10628
rect 14461 10619 14519 10625
rect 14660 10600 14688 10628
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 15102 10656 15108 10668
rect 14936 10628 15108 10656
rect 12584 10560 13584 10588
rect 13924 10560 14412 10588
rect 12584 10548 12590 10560
rect 7926 10520 7932 10532
rect 6380 10492 7932 10520
rect 7926 10480 7932 10492
rect 7984 10480 7990 10532
rect 11238 10520 11244 10532
rect 8312 10492 11244 10520
rect 992 10424 3648 10452
rect 4801 10455 4859 10461
rect 992 10412 998 10424
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 4890 10452 4896 10464
rect 4847 10424 4896 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 6196 10452 6224 10480
rect 8312 10452 8340 10492
rect 11238 10480 11244 10492
rect 11296 10480 11302 10532
rect 13357 10523 13415 10529
rect 13357 10489 13369 10523
rect 13403 10520 13415 10523
rect 13446 10520 13452 10532
rect 13403 10492 13452 10520
rect 13403 10489 13415 10492
rect 13357 10483 13415 10489
rect 13446 10480 13452 10492
rect 13504 10480 13510 10532
rect 13556 10520 13584 10560
rect 14642 10548 14648 10600
rect 14700 10548 14706 10600
rect 14936 10520 14964 10628
rect 15102 10616 15108 10628
rect 15160 10656 15166 10668
rect 15657 10659 15715 10665
rect 15657 10656 15669 10659
rect 15160 10628 15669 10656
rect 15160 10616 15166 10628
rect 15657 10625 15669 10628
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 15010 10548 15016 10600
rect 15068 10588 15074 10600
rect 15948 10588 15976 10619
rect 15068 10560 15976 10588
rect 15068 10548 15074 10560
rect 15470 10520 15476 10532
rect 13556 10492 14964 10520
rect 15431 10492 15476 10520
rect 15470 10480 15476 10492
rect 15528 10480 15534 10532
rect 15654 10480 15660 10532
rect 15712 10520 15718 10532
rect 16040 10520 16068 10696
rect 15712 10492 16068 10520
rect 15712 10480 15718 10492
rect 6196 10424 8340 10452
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 8570 10452 8576 10464
rect 8444 10424 8576 10452
rect 8444 10412 8450 10424
rect 8570 10412 8576 10424
rect 8628 10452 8634 10464
rect 9125 10455 9183 10461
rect 9125 10452 9137 10455
rect 8628 10424 9137 10452
rect 8628 10412 8634 10424
rect 9125 10421 9137 10424
rect 9171 10421 9183 10455
rect 9125 10415 9183 10421
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 10502 10452 10508 10464
rect 10192 10424 10508 10452
rect 10192 10412 10198 10424
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 10778 10412 10784 10464
rect 10836 10452 10842 10464
rect 12250 10452 12256 10464
rect 10836 10424 12256 10452
rect 10836 10412 10842 10424
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 13170 10452 13176 10464
rect 12492 10424 13176 10452
rect 12492 10412 12498 10424
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 14090 10452 14096 10464
rect 13596 10424 14096 10452
rect 13596 10412 13602 10424
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 16850 10452 16856 10464
rect 14240 10424 16856 10452
rect 14240 10412 14246 10424
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 1104 10362 16836 10384
rect 1104 10310 2924 10362
rect 2976 10310 2988 10362
rect 3040 10310 3052 10362
rect 3104 10310 3116 10362
rect 3168 10310 3180 10362
rect 3232 10310 6872 10362
rect 6924 10310 6936 10362
rect 6988 10310 7000 10362
rect 7052 10310 7064 10362
rect 7116 10310 7128 10362
rect 7180 10310 10820 10362
rect 10872 10310 10884 10362
rect 10936 10310 10948 10362
rect 11000 10310 11012 10362
rect 11064 10310 11076 10362
rect 11128 10310 14768 10362
rect 14820 10310 14832 10362
rect 14884 10310 14896 10362
rect 14948 10310 14960 10362
rect 15012 10310 15024 10362
rect 15076 10310 16836 10362
rect 1104 10288 16836 10310
rect 3878 10248 3884 10260
rect 3839 10220 3884 10248
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 5166 10248 5172 10260
rect 4540 10220 5172 10248
rect 1394 10180 1400 10192
rect 1320 10152 1400 10180
rect 1320 9976 1348 10152
rect 1394 10140 1400 10152
rect 1452 10140 1458 10192
rect 4540 10180 4568 10220
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 8110 10248 8116 10260
rect 8071 10220 8116 10248
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 11330 10248 11336 10260
rect 9364 10220 11336 10248
rect 9364 10208 9370 10220
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 11701 10251 11759 10257
rect 11701 10248 11713 10251
rect 11572 10220 11713 10248
rect 11572 10208 11578 10220
rect 11701 10217 11713 10220
rect 11747 10217 11759 10251
rect 11701 10211 11759 10217
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 12032 10220 12472 10248
rect 12032 10208 12038 10220
rect 3252 10152 4568 10180
rect 1486 10112 1492 10124
rect 1447 10084 1492 10112
rect 1486 10072 1492 10084
rect 1544 10072 1550 10124
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 3252 10121 3280 10152
rect 5718 10140 5724 10192
rect 5776 10180 5782 10192
rect 5902 10180 5908 10192
rect 5776 10152 5908 10180
rect 5776 10140 5782 10152
rect 5902 10140 5908 10152
rect 5960 10140 5966 10192
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 8294 10180 8300 10192
rect 6236 10152 8300 10180
rect 6236 10140 6242 10152
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 9950 10140 9956 10192
rect 10008 10180 10014 10192
rect 12444 10180 12472 10220
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13906 10248 13912 10260
rect 12860 10220 13912 10248
rect 12860 10208 12866 10220
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 14016 10220 14688 10248
rect 14016 10180 14044 10220
rect 10008 10152 12388 10180
rect 12444 10152 14044 10180
rect 10008 10140 10014 10152
rect 3237 10115 3295 10121
rect 3237 10112 3249 10115
rect 3200 10084 3249 10112
rect 3200 10072 3206 10084
rect 3237 10081 3249 10084
rect 3283 10081 3295 10115
rect 3237 10075 3295 10081
rect 4062 10072 4068 10124
rect 4120 10112 4126 10124
rect 4709 10115 4767 10121
rect 4709 10112 4721 10115
rect 4120 10084 4721 10112
rect 4120 10072 4126 10084
rect 4709 10081 4721 10084
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 9030 10112 9036 10124
rect 5132 10084 9036 10112
rect 5132 10072 5138 10084
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 9401 10115 9459 10121
rect 9401 10081 9413 10115
rect 9447 10112 9459 10115
rect 12360 10112 12388 10152
rect 14090 10140 14096 10192
rect 14148 10180 14154 10192
rect 14550 10180 14556 10192
rect 14148 10152 14556 10180
rect 14148 10140 14154 10152
rect 14550 10140 14556 10152
rect 14608 10140 14614 10192
rect 14660 10180 14688 10220
rect 14734 10208 14740 10260
rect 14792 10248 14798 10260
rect 15470 10248 15476 10260
rect 14792 10220 15476 10248
rect 14792 10208 14798 10220
rect 15470 10208 15476 10220
rect 15528 10208 15534 10260
rect 15654 10208 15660 10260
rect 15712 10248 15718 10260
rect 16390 10248 16396 10260
rect 15712 10220 16396 10248
rect 15712 10208 15718 10220
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 15749 10183 15807 10189
rect 15749 10180 15761 10183
rect 14660 10152 15761 10180
rect 15749 10149 15761 10152
rect 15795 10149 15807 10183
rect 15749 10143 15807 10149
rect 13262 10112 13268 10124
rect 9447 10084 12296 10112
rect 12360 10084 13268 10112
rect 9447 10081 9459 10084
rect 9401 10075 9459 10081
rect 3694 10004 3700 10056
rect 3752 10044 3758 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3752 10016 3801 10044
rect 3752 10004 3758 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 1765 9979 1823 9985
rect 1765 9976 1777 9979
rect 1320 9948 1777 9976
rect 1765 9945 1777 9948
rect 1811 9945 1823 9979
rect 1765 9939 1823 9945
rect 1780 9908 1808 9939
rect 2774 9936 2780 9988
rect 2832 9936 2838 9988
rect 3326 9936 3332 9988
rect 3384 9976 3390 9988
rect 3988 9976 4016 10007
rect 4246 10004 4252 10056
rect 4304 10044 4310 10056
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 4304 10016 4445 10044
rect 4304 10004 4310 10016
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 6730 10044 6736 10056
rect 6687 10016 6736 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 6730 10004 6736 10016
rect 6788 10044 6794 10056
rect 7190 10044 7196 10056
rect 6788 10016 7196 10044
rect 6788 10004 6794 10016
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8754 10044 8760 10056
rect 7984 10016 8760 10044
rect 7984 10004 7990 10016
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 11422 10044 11428 10056
rect 9171 10016 11428 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 11422 10004 11428 10016
rect 11480 10044 11486 10056
rect 12066 10044 12072 10056
rect 11480 10016 12072 10044
rect 11480 10004 11486 10016
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12268 10044 12296 10084
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 14568 10112 14596 10140
rect 14568 10084 14780 10112
rect 12526 10044 12532 10056
rect 12268 10016 12532 10044
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10044 12771 10047
rect 12802 10044 12808 10056
rect 12759 10016 12808 10044
rect 12759 10013 12771 10016
rect 12713 10007 12771 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 12986 10044 12992 10056
rect 12947 10016 12992 10044
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 14550 10044 14556 10056
rect 13096 10016 14136 10044
rect 14511 10016 14556 10044
rect 6086 9976 6092 9988
rect 3384 9948 4016 9976
rect 5934 9948 6092 9976
rect 3384 9936 3390 9948
rect 6086 9936 6092 9948
rect 6144 9936 6150 9988
rect 10413 9979 10471 9985
rect 10413 9945 10425 9979
rect 10459 9976 10471 9979
rect 10502 9976 10508 9988
rect 10459 9948 10508 9976
rect 10459 9945 10471 9948
rect 10413 9939 10471 9945
rect 10502 9936 10508 9948
rect 10560 9936 10566 9988
rect 13096 9976 13124 10016
rect 11256 9948 13124 9976
rect 4154 9908 4160 9920
rect 1780 9880 4160 9908
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 6181 9911 6239 9917
rect 6181 9877 6193 9911
rect 6227 9908 6239 9911
rect 6362 9908 6368 9920
rect 6227 9880 6368 9908
rect 6227 9877 6239 9880
rect 6181 9871 6239 9877
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 8570 9868 8576 9920
rect 8628 9908 8634 9920
rect 11256 9908 11284 9948
rect 13630 9936 13636 9988
rect 13688 9976 13694 9988
rect 13814 9976 13820 9988
rect 13688 9948 13820 9976
rect 13688 9936 13694 9948
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 14108 9976 14136 10016
rect 14550 10004 14556 10016
rect 14608 10004 14614 10056
rect 14752 10053 14780 10084
rect 15470 10072 15476 10124
rect 15528 10112 15534 10124
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 15528 10084 15669 10112
rect 15528 10072 15534 10084
rect 15657 10081 15669 10084
rect 15703 10112 15715 10115
rect 16206 10112 16212 10124
rect 15703 10084 16212 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 14918 10053 14924 10056
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10013 14795 10047
rect 14737 10007 14795 10013
rect 14901 10047 14924 10053
rect 14901 10013 14913 10047
rect 14901 10007 14924 10013
rect 14918 10004 14924 10007
rect 14976 10004 14982 10056
rect 15565 10047 15623 10053
rect 15565 10013 15577 10047
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10044 15899 10047
rect 16850 10044 16856 10056
rect 15887 10016 16856 10044
rect 15887 10013 15899 10016
rect 15841 10007 15899 10013
rect 14645 9979 14703 9985
rect 14645 9976 14657 9979
rect 14108 9948 14657 9976
rect 14645 9945 14657 9948
rect 14691 9976 14703 9979
rect 15197 9979 15255 9985
rect 15197 9976 15209 9979
rect 14691 9948 15209 9976
rect 14691 9945 14703 9948
rect 14645 9939 14703 9945
rect 15197 9945 15209 9948
rect 15243 9945 15255 9979
rect 15580 9976 15608 10007
rect 16850 10004 16856 10016
rect 16908 10004 16914 10056
rect 15746 9976 15752 9988
rect 15580 9948 15752 9976
rect 15197 9939 15255 9945
rect 15746 9936 15752 9948
rect 15804 9976 15810 9988
rect 16390 9976 16396 9988
rect 15804 9948 16396 9976
rect 15804 9936 15810 9948
rect 16390 9936 16396 9948
rect 16448 9936 16454 9988
rect 8628 9880 11284 9908
rect 8628 9868 8634 9880
rect 11422 9868 11428 9920
rect 11480 9908 11486 9920
rect 14274 9908 14280 9920
rect 11480 9880 14280 9908
rect 11480 9868 11486 9880
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 14366 9868 14372 9920
rect 14424 9908 14430 9920
rect 14424 9880 14469 9908
rect 14424 9868 14430 9880
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 15381 9911 15439 9917
rect 15381 9908 15393 9911
rect 14608 9880 15393 9908
rect 14608 9868 14614 9880
rect 15381 9877 15393 9880
rect 15427 9877 15439 9911
rect 15381 9871 15439 9877
rect 1104 9818 16836 9840
rect 1104 9766 4898 9818
rect 4950 9766 4962 9818
rect 5014 9766 5026 9818
rect 5078 9766 5090 9818
rect 5142 9766 5154 9818
rect 5206 9766 8846 9818
rect 8898 9766 8910 9818
rect 8962 9766 8974 9818
rect 9026 9766 9038 9818
rect 9090 9766 9102 9818
rect 9154 9766 12794 9818
rect 12846 9766 12858 9818
rect 12910 9766 12922 9818
rect 12974 9766 12986 9818
rect 13038 9766 13050 9818
rect 13102 9766 16836 9818
rect 1104 9744 16836 9766
rect 1026 9664 1032 9716
rect 1084 9704 1090 9716
rect 1578 9704 1584 9716
rect 1084 9676 1584 9704
rect 1084 9664 1090 9676
rect 1578 9664 1584 9676
rect 1636 9664 1642 9716
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 9582 9704 9588 9716
rect 4120 9676 9588 9704
rect 4120 9664 4126 9676
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 10318 9664 10324 9716
rect 10376 9704 10382 9716
rect 10594 9704 10600 9716
rect 10376 9676 10600 9704
rect 10376 9664 10382 9676
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 11330 9664 11336 9716
rect 11388 9704 11394 9716
rect 11388 9676 12848 9704
rect 11388 9664 11394 9676
rect 2314 9596 2320 9648
rect 2372 9636 2378 9648
rect 5902 9636 5908 9648
rect 2372 9608 4108 9636
rect 2372 9596 2378 9608
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3234 9568 3240 9580
rect 3007 9540 3240 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 4080 9577 4108 9608
rect 5092 9608 5908 9636
rect 5092 9577 5120 9608
rect 5902 9596 5908 9608
rect 5960 9596 5966 9648
rect 7282 9636 7288 9648
rect 6564 9608 7288 9636
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5442 9568 5448 9580
rect 5077 9531 5135 9537
rect 5184 9540 5448 9568
rect 2041 9503 2099 9509
rect 2041 9469 2053 9503
rect 2087 9500 2099 9503
rect 2130 9500 2136 9512
rect 2087 9472 2136 9500
rect 2087 9469 2099 9472
rect 2041 9463 2099 9469
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2593 9503 2651 9509
rect 2593 9500 2605 9503
rect 2363 9472 2605 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2593 9469 2605 9472
rect 2639 9500 2651 9503
rect 3142 9500 3148 9512
rect 2639 9472 3148 9500
rect 2639 9469 2651 9472
rect 2593 9463 2651 9469
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 2774 9392 2780 9444
rect 2832 9432 2838 9444
rect 2869 9435 2927 9441
rect 2869 9432 2881 9435
rect 2832 9404 2881 9432
rect 2832 9392 2838 9404
rect 2869 9401 2881 9404
rect 2915 9401 2927 9435
rect 2869 9395 2927 9401
rect 3712 9364 3740 9531
rect 3789 9503 3847 9509
rect 3789 9469 3801 9503
rect 3835 9469 3847 9503
rect 3789 9463 3847 9469
rect 3804 9432 3832 9463
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3936 9472 3985 9500
rect 3936 9460 3942 9472
rect 3973 9469 3985 9472
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 5184 9432 5212 9540
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 6564 9577 6592 9608
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 8846 9636 8852 9648
rect 8168 9608 8852 9636
rect 8168 9596 8174 9608
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 9217 9639 9275 9645
rect 9217 9605 9229 9639
rect 9263 9636 9275 9639
rect 11974 9636 11980 9648
rect 9263 9608 11980 9636
rect 9263 9605 9275 9608
rect 9217 9599 9275 9605
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 6549 9571 6607 9577
rect 6288 9540 6500 9568
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 6086 9500 6092 9512
rect 5399 9472 6092 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 6086 9460 6092 9472
rect 6144 9460 6150 9512
rect 3804 9404 5212 9432
rect 5261 9435 5319 9441
rect 5261 9401 5273 9435
rect 5307 9432 5319 9435
rect 6288 9432 6316 9540
rect 6362 9460 6368 9512
rect 6420 9460 6426 9512
rect 6472 9500 6500 9540
rect 6549 9537 6561 9571
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9568 7067 9571
rect 11238 9568 11244 9580
rect 7055 9540 11244 9568
rect 7055 9537 7067 9540
rect 7009 9531 7067 9537
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9568 11575 9571
rect 11606 9568 11612 9580
rect 11563 9540 11612 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 11784 9571 11842 9577
rect 11784 9537 11796 9571
rect 11830 9568 11842 9571
rect 12342 9568 12348 9580
rect 11830 9540 12348 9568
rect 11830 9537 11842 9540
rect 11784 9531 11842 9537
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 12820 9568 12848 9676
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 14737 9707 14795 9713
rect 13320 9676 13860 9704
rect 13320 9664 13326 9676
rect 12894 9596 12900 9648
rect 12952 9636 12958 9648
rect 13832 9636 13860 9676
rect 14737 9673 14749 9707
rect 14783 9704 14795 9707
rect 14826 9704 14832 9716
rect 14783 9676 14832 9704
rect 14783 9673 14795 9676
rect 14737 9667 14795 9673
rect 14826 9664 14832 9676
rect 14884 9664 14890 9716
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 15930 9704 15936 9716
rect 15344 9676 15936 9704
rect 15344 9664 15350 9676
rect 15930 9664 15936 9676
rect 15988 9664 15994 9716
rect 12952 9608 13768 9636
rect 13832 9608 15424 9636
rect 12952 9596 12958 9608
rect 13613 9571 13671 9577
rect 13613 9568 13625 9571
rect 12820 9540 13625 9568
rect 13613 9537 13625 9540
rect 13659 9537 13671 9571
rect 13740 9568 13768 9608
rect 15194 9568 15200 9580
rect 13740 9540 15200 9568
rect 13613 9531 13671 9537
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15396 9577 15424 9608
rect 15381 9571 15439 9577
rect 15381 9537 15393 9571
rect 15427 9537 15439 9571
rect 15381 9531 15439 9537
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 9950 9500 9956 9512
rect 6472 9472 9956 9500
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 10978 9460 10984 9512
rect 11036 9500 11042 9512
rect 11330 9500 11336 9512
rect 11036 9472 11336 9500
rect 11036 9460 11042 9472
rect 11330 9460 11336 9472
rect 11388 9460 11394 9512
rect 13354 9500 13360 9512
rect 13315 9472 13360 9500
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 5307 9404 6316 9432
rect 6380 9432 6408 9460
rect 8297 9435 8355 9441
rect 8297 9432 8309 9435
rect 6380 9404 8309 9432
rect 5307 9401 5319 9404
rect 5261 9395 5319 9401
rect 8297 9401 8309 9404
rect 8343 9401 8355 9435
rect 8297 9395 8355 9401
rect 9398 9392 9404 9444
rect 9456 9432 9462 9444
rect 11514 9432 11520 9444
rect 9456 9404 11520 9432
rect 9456 9392 9462 9404
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 12526 9392 12532 9444
rect 12584 9432 12590 9444
rect 12894 9432 12900 9444
rect 12584 9404 12900 9432
rect 12584 9392 12590 9404
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 15580 9432 15608 9531
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 15712 9540 15757 9568
rect 15712 9528 15718 9540
rect 14292 9404 15608 9432
rect 4154 9364 4160 9376
rect 3712 9336 4160 9364
rect 4154 9324 4160 9336
rect 4212 9364 4218 9376
rect 4798 9364 4804 9376
rect 4212 9336 4804 9364
rect 4212 9324 4218 9336
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5442 9364 5448 9376
rect 5215 9336 5448 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 6822 9364 6828 9376
rect 6411 9336 6828 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 10502 9364 10508 9376
rect 8720 9336 10508 9364
rect 8720 9324 8726 9336
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 10594 9324 10600 9376
rect 10652 9364 10658 9376
rect 14292 9364 14320 9404
rect 10652 9336 14320 9364
rect 15197 9367 15255 9373
rect 10652 9324 10658 9336
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 15654 9364 15660 9376
rect 15243 9336 15660 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 1104 9274 16836 9296
rect 1104 9222 2924 9274
rect 2976 9222 2988 9274
rect 3040 9222 3052 9274
rect 3104 9222 3116 9274
rect 3168 9222 3180 9274
rect 3232 9222 6872 9274
rect 6924 9222 6936 9274
rect 6988 9222 7000 9274
rect 7052 9222 7064 9274
rect 7116 9222 7128 9274
rect 7180 9222 10820 9274
rect 10872 9222 10884 9274
rect 10936 9222 10948 9274
rect 11000 9222 11012 9274
rect 11064 9222 11076 9274
rect 11128 9222 14768 9274
rect 14820 9222 14832 9274
rect 14884 9222 14896 9274
rect 14948 9222 14960 9274
rect 15012 9222 15024 9274
rect 15076 9222 16836 9274
rect 1104 9200 16836 9222
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 6086 9160 6092 9172
rect 3283 9132 6092 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 6270 9160 6276 9172
rect 6231 9132 6276 9160
rect 6270 9120 6276 9132
rect 6328 9120 6334 9172
rect 7926 9160 7932 9172
rect 6656 9132 7932 9160
rect 6656 9092 6684 9132
rect 7926 9120 7932 9132
rect 7984 9160 7990 9172
rect 8389 9163 8447 9169
rect 8389 9160 8401 9163
rect 7984 9132 8401 9160
rect 7984 9120 7990 9132
rect 8389 9129 8401 9132
rect 8435 9129 8447 9163
rect 8389 9123 8447 9129
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 14093 9163 14151 9169
rect 14093 9160 14105 9163
rect 8628 9132 14105 9160
rect 8628 9120 8634 9132
rect 14093 9129 14105 9132
rect 14139 9129 14151 9163
rect 15562 9160 15568 9172
rect 14093 9123 14151 9129
rect 14384 9132 15568 9160
rect 3804 9064 6684 9092
rect 1489 9027 1547 9033
rect 1489 8993 1501 9027
rect 1535 9024 1547 9027
rect 2130 9024 2136 9036
rect 1535 8996 2136 9024
rect 1535 8993 1547 8996
rect 1489 8987 1547 8993
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 3804 8965 3832 9064
rect 9214 9052 9220 9104
rect 9272 9092 9278 9104
rect 10594 9092 10600 9104
rect 9272 9064 10600 9092
rect 9272 9052 9278 9064
rect 10594 9052 10600 9064
rect 10652 9052 10658 9104
rect 11330 9092 11336 9104
rect 10704 9064 11336 9092
rect 4430 9024 4436 9036
rect 3988 8996 4436 9024
rect 3988 8965 4016 8996
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 5810 9024 5816 9036
rect 4724 8996 5816 9024
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4724 8956 4752 8996
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 6546 8984 6552 9036
rect 6604 9024 6610 9036
rect 7009 9027 7067 9033
rect 7009 9024 7021 9027
rect 6604 8996 7021 9024
rect 6604 8984 6610 8996
rect 7009 8993 7021 8996
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 8846 8984 8852 9036
rect 8904 9024 8910 9036
rect 8904 8996 9444 9024
rect 8904 8984 8910 8996
rect 4203 8928 4752 8956
rect 4801 8959 4859 8965
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4801 8925 4813 8959
rect 4847 8956 4859 8959
rect 6730 8956 6736 8968
rect 4847 8928 6736 8956
rect 4847 8925 4859 8928
rect 4801 8919 4859 8925
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 7156 8928 7604 8956
rect 7156 8916 7162 8928
rect 1026 8848 1032 8900
rect 1084 8888 1090 8900
rect 1765 8891 1823 8897
rect 1765 8888 1777 8891
rect 1084 8860 1777 8888
rect 1084 8848 1090 8860
rect 1765 8857 1777 8860
rect 1811 8857 1823 8891
rect 3878 8888 3884 8900
rect 2990 8860 3884 8888
rect 1765 8851 1823 8857
rect 3878 8848 3884 8860
rect 3936 8848 3942 8900
rect 4065 8891 4123 8897
rect 4065 8857 4077 8891
rect 4111 8888 4123 8891
rect 6638 8888 6644 8900
rect 4111 8860 6644 8888
rect 4111 8857 4123 8860
rect 4065 8851 4123 8857
rect 6638 8848 6644 8860
rect 6696 8848 6702 8900
rect 7276 8891 7334 8897
rect 7276 8857 7288 8891
rect 7322 8888 7334 8891
rect 7466 8888 7472 8900
rect 7322 8860 7472 8888
rect 7322 8857 7334 8860
rect 7276 8851 7334 8857
rect 7466 8848 7472 8860
rect 7524 8848 7530 8900
rect 7576 8888 7604 8928
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 7800 8928 9321 8956
rect 7800 8916 7806 8928
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9416 8956 9444 8996
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 10704 9024 10732 9064
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 12526 9052 12532 9104
rect 12584 9092 12590 9104
rect 12802 9092 12808 9104
rect 12584 9064 12808 9092
rect 12584 9052 12590 9064
rect 12802 9052 12808 9064
rect 12860 9092 12866 9104
rect 12860 9064 14136 9092
rect 12860 9052 12866 9064
rect 14108 9036 14136 9064
rect 9640 8996 10732 9024
rect 9640 8984 9646 8996
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11517 9027 11575 9033
rect 11517 9024 11529 9027
rect 11204 8996 11529 9024
rect 11204 8984 11210 8996
rect 11517 8993 11529 8996
rect 11563 8993 11575 9027
rect 11517 8987 11575 8993
rect 12710 8984 12716 9036
rect 12768 9024 12774 9036
rect 12768 8996 13400 9024
rect 12768 8984 12774 8996
rect 12986 8956 12992 8968
rect 9416 8928 12992 8956
rect 9309 8919 9367 8925
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 13372 8965 13400 8996
rect 14090 8984 14096 9036
rect 14148 8984 14154 9036
rect 14274 9024 14280 9036
rect 14235 8996 14280 9024
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 14384 9033 14412 9132
rect 15562 9120 15568 9132
rect 15620 9120 15626 9172
rect 15930 9092 15936 9104
rect 14476 9064 15936 9092
rect 14476 9033 14504 9064
rect 15930 9052 15936 9064
rect 15988 9052 15994 9104
rect 14369 9027 14427 9033
rect 14369 8993 14381 9027
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 14461 9027 14519 9033
rect 14461 8993 14473 9027
rect 14507 8993 14519 9027
rect 14461 8987 14519 8993
rect 14826 8984 14832 9036
rect 14884 9024 14890 9036
rect 14884 8996 15332 9024
rect 14884 8984 14890 8996
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 13722 8956 13728 8968
rect 13495 8928 13728 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 14553 8959 14611 8965
rect 14553 8956 14565 8959
rect 14056 8928 14565 8956
rect 14056 8916 14062 8928
rect 14553 8925 14565 8928
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 14642 8916 14648 8968
rect 14700 8956 14706 8968
rect 15010 8956 15016 8968
rect 14700 8928 15016 8956
rect 14700 8916 14706 8928
rect 15010 8916 15016 8928
rect 15068 8956 15074 8968
rect 15304 8965 15332 8996
rect 15289 8959 15347 8965
rect 15068 8928 15240 8956
rect 15068 8916 15074 8928
rect 7576 8860 10916 8888
rect 4338 8820 4344 8832
rect 4299 8792 4344 8820
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 6086 8780 6092 8832
rect 6144 8820 6150 8832
rect 9306 8820 9312 8832
rect 6144 8792 9312 8820
rect 6144 8780 6150 8792
rect 9306 8780 9312 8792
rect 9364 8780 9370 8832
rect 10778 8820 10784 8832
rect 10739 8792 10784 8820
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 10888 8820 10916 8860
rect 11146 8848 11152 8900
rect 11204 8888 11210 8900
rect 11422 8888 11428 8900
rect 11204 8860 11428 8888
rect 11204 8848 11210 8860
rect 11422 8848 11428 8860
rect 11480 8848 11486 8900
rect 11784 8891 11842 8897
rect 11784 8857 11796 8891
rect 11830 8888 11842 8891
rect 11974 8888 11980 8900
rect 11830 8860 11980 8888
rect 11830 8857 11842 8860
rect 11784 8851 11842 8857
rect 11974 8848 11980 8860
rect 12032 8848 12038 8900
rect 12342 8848 12348 8900
rect 12400 8888 12406 8900
rect 15105 8891 15163 8897
rect 15105 8888 15117 8891
rect 12400 8860 15117 8888
rect 12400 8848 12406 8860
rect 15105 8857 15117 8860
rect 15151 8857 15163 8891
rect 15212 8888 15240 8928
rect 15289 8925 15301 8959
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 15565 8959 15623 8965
rect 15565 8925 15577 8959
rect 15611 8956 15623 8959
rect 15746 8956 15752 8968
rect 15611 8928 15752 8956
rect 15611 8925 15623 8928
rect 15565 8919 15623 8925
rect 15746 8916 15752 8928
rect 15804 8956 15810 8968
rect 16206 8956 16212 8968
rect 15804 8928 16212 8956
rect 15804 8916 15810 8928
rect 16206 8916 16212 8928
rect 16264 8916 16270 8968
rect 15473 8891 15531 8897
rect 15473 8888 15485 8891
rect 15212 8860 15485 8888
rect 15105 8851 15163 8857
rect 15473 8857 15485 8860
rect 15519 8857 15531 8891
rect 15473 8851 15531 8857
rect 12897 8823 12955 8829
rect 12897 8820 12909 8823
rect 10888 8792 12909 8820
rect 12897 8789 12909 8792
rect 12943 8820 12955 8823
rect 15378 8820 15384 8832
rect 12943 8792 15384 8820
rect 12943 8789 12955 8792
rect 12897 8783 12955 8789
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 1104 8730 16836 8752
rect 1104 8678 4898 8730
rect 4950 8678 4962 8730
rect 5014 8678 5026 8730
rect 5078 8678 5090 8730
rect 5142 8678 5154 8730
rect 5206 8678 8846 8730
rect 8898 8678 8910 8730
rect 8962 8678 8974 8730
rect 9026 8678 9038 8730
rect 9090 8678 9102 8730
rect 9154 8678 12794 8730
rect 12846 8678 12858 8730
rect 12910 8678 12922 8730
rect 12974 8678 12986 8730
rect 13038 8678 13050 8730
rect 13102 8678 16836 8730
rect 1104 8656 16836 8678
rect 3329 8619 3387 8625
rect 3329 8585 3341 8619
rect 3375 8616 3387 8619
rect 3602 8616 3608 8628
rect 3375 8588 3608 8616
rect 3375 8585 3387 8588
rect 3329 8579 3387 8585
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 9582 8616 9588 8628
rect 4448 8588 9588 8616
rect 4448 8548 4476 8588
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 12434 8616 12440 8628
rect 10784 8588 12440 8616
rect 3082 8520 4476 8548
rect 5442 8508 5448 8560
rect 5500 8548 5506 8560
rect 6362 8548 6368 8560
rect 5500 8520 6368 8548
rect 5500 8508 5506 8520
rect 6362 8508 6368 8520
rect 6420 8508 6426 8560
rect 10784 8548 10812 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13446 8616 13452 8628
rect 13403 8588 13452 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 13538 8576 13544 8628
rect 13596 8576 13602 8628
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 15197 8619 15255 8625
rect 15197 8616 15209 8619
rect 14792 8588 15209 8616
rect 14792 8576 14798 8588
rect 15197 8585 15209 8588
rect 15243 8585 15255 8619
rect 15197 8579 15255 8585
rect 7866 8520 10812 8548
rect 10870 8508 10876 8560
rect 10928 8548 10934 8560
rect 12894 8548 12900 8560
rect 10928 8520 12900 8548
rect 10928 8508 10934 8520
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 3789 8483 3847 8489
rect 3789 8480 3801 8483
rect 3660 8452 3801 8480
rect 3660 8440 3666 8452
rect 3789 8449 3801 8452
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 5166 8440 5172 8492
rect 5224 8440 5230 8492
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8352 8452 8861 8480
rect 8352 8440 8358 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 10410 8480 10416 8492
rect 10371 8452 10416 8480
rect 8849 8443 8907 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 10520 8452 11529 8480
rect 1578 8412 1584 8424
rect 1539 8384 1584 8412
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 4062 8412 4068 8424
rect 1903 8384 3740 8412
rect 4023 8384 4068 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 2038 8236 2044 8288
rect 2096 8276 2102 8288
rect 2314 8276 2320 8288
rect 2096 8248 2320 8276
rect 2096 8236 2102 8248
rect 2314 8236 2320 8248
rect 2372 8236 2378 8288
rect 3712 8285 3740 8384
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4430 8372 4436 8424
rect 4488 8412 4494 8424
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 4488 8384 5549 8412
rect 4488 8372 4494 8384
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 6362 8412 6368 8424
rect 6323 8384 6368 8412
rect 5537 8375 5595 8381
rect 6362 8372 6368 8384
rect 6420 8372 6426 8424
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 6687 8384 9536 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 5074 8304 5080 8356
rect 5132 8344 5138 8356
rect 9508 8344 9536 8384
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 10520 8412 10548 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11784 8483 11842 8489
rect 11784 8449 11796 8483
rect 11830 8480 11842 8483
rect 12342 8480 12348 8492
rect 11830 8452 12348 8480
rect 11830 8449 11842 8452
rect 11784 8443 11842 8449
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 12802 8440 12808 8492
rect 12860 8480 12866 8492
rect 13556 8480 13584 8576
rect 13722 8548 13728 8560
rect 13683 8520 13728 8548
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 14642 8508 14648 8560
rect 14700 8548 14706 8560
rect 15212 8548 15240 8579
rect 14700 8520 15148 8548
rect 15212 8520 15700 8548
rect 14700 8508 14706 8520
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 12860 8452 13584 8480
rect 14200 8452 14565 8480
rect 12860 8440 12866 8452
rect 9640 8384 10548 8412
rect 9640 8372 9646 8384
rect 11330 8372 11336 8424
rect 11388 8372 11394 8424
rect 13817 8415 13875 8421
rect 13817 8412 13829 8415
rect 12544 8384 13829 8412
rect 11348 8344 11376 8372
rect 5132 8316 6224 8344
rect 5132 8304 5138 8316
rect 3697 8279 3755 8285
rect 3697 8245 3709 8279
rect 3743 8276 3755 8279
rect 6086 8276 6092 8288
rect 3743 8248 6092 8276
rect 3743 8245 3755 8248
rect 3697 8239 3755 8245
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 6196 8276 6224 8316
rect 7659 8316 8432 8344
rect 9508 8316 11376 8344
rect 7659 8276 7687 8316
rect 6196 8248 7687 8276
rect 8113 8279 8171 8285
rect 8113 8245 8125 8279
rect 8159 8276 8171 8279
rect 8294 8276 8300 8288
rect 8159 8248 8300 8276
rect 8159 8245 8171 8248
rect 8113 8239 8171 8245
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 8404 8276 8432 8316
rect 11330 8276 11336 8288
rect 8404 8248 11336 8276
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11514 8236 11520 8288
rect 11572 8276 11578 8288
rect 12544 8276 12572 8384
rect 13817 8381 13829 8384
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8412 14059 8415
rect 14090 8412 14096 8424
rect 14047 8384 14096 8412
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 13078 8304 13084 8356
rect 13136 8344 13142 8356
rect 13538 8344 13544 8356
rect 13136 8316 13544 8344
rect 13136 8304 13142 8316
rect 13538 8304 13544 8316
rect 13596 8304 13602 8356
rect 13630 8304 13636 8356
rect 13688 8344 13694 8356
rect 14200 8344 14228 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 15120 8480 15148 8520
rect 15565 8483 15623 8489
rect 15565 8480 15577 8483
rect 15120 8452 15577 8480
rect 14553 8443 14611 8449
rect 15565 8449 15577 8452
rect 15611 8449 15623 8483
rect 15565 8443 15623 8449
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8412 14703 8415
rect 14734 8412 14740 8424
rect 14691 8384 14740 8412
rect 14691 8381 14703 8384
rect 14645 8375 14703 8381
rect 14734 8372 14740 8384
rect 14792 8372 14798 8424
rect 15672 8421 15700 8520
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 16390 8480 16396 8492
rect 15887 8452 16396 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16390 8440 16396 8452
rect 16448 8440 16454 8492
rect 15657 8415 15715 8421
rect 15657 8381 15669 8415
rect 15703 8381 15715 8415
rect 15657 8375 15715 8381
rect 15746 8372 15752 8424
rect 15804 8372 15810 8424
rect 13688 8316 14228 8344
rect 14921 8347 14979 8353
rect 13688 8304 13694 8316
rect 14921 8313 14933 8347
rect 14967 8344 14979 8347
rect 15102 8344 15108 8356
rect 14967 8316 15108 8344
rect 14967 8313 14979 8316
rect 14921 8307 14979 8313
rect 15102 8304 15108 8316
rect 15160 8304 15166 8356
rect 15286 8304 15292 8356
rect 15344 8344 15350 8356
rect 15764 8344 15792 8372
rect 15344 8316 15792 8344
rect 15344 8304 15350 8316
rect 11572 8248 12572 8276
rect 12897 8279 12955 8285
rect 11572 8236 11578 8248
rect 12897 8245 12909 8279
rect 12943 8276 12955 8279
rect 15010 8276 15016 8288
rect 12943 8248 15016 8276
rect 12943 8245 12955 8248
rect 12897 8239 12955 8245
rect 15010 8236 15016 8248
rect 15068 8236 15074 8288
rect 15565 8279 15623 8285
rect 15565 8245 15577 8279
rect 15611 8276 15623 8279
rect 15672 8276 15700 8316
rect 15611 8248 15700 8276
rect 16025 8279 16083 8285
rect 15611 8245 15623 8248
rect 15565 8239 15623 8245
rect 16025 8245 16037 8279
rect 16071 8276 16083 8279
rect 17678 8276 17684 8288
rect 16071 8248 17684 8276
rect 16071 8245 16083 8248
rect 16025 8239 16083 8245
rect 17678 8236 17684 8248
rect 17736 8236 17742 8288
rect 1104 8186 16836 8208
rect 1104 8134 2924 8186
rect 2976 8134 2988 8186
rect 3040 8134 3052 8186
rect 3104 8134 3116 8186
rect 3168 8134 3180 8186
rect 3232 8134 6872 8186
rect 6924 8134 6936 8186
rect 6988 8134 7000 8186
rect 7052 8134 7064 8186
rect 7116 8134 7128 8186
rect 7180 8134 10820 8186
rect 10872 8134 10884 8186
rect 10936 8134 10948 8186
rect 11000 8134 11012 8186
rect 11064 8134 11076 8186
rect 11128 8134 14768 8186
rect 14820 8134 14832 8186
rect 14884 8134 14896 8186
rect 14948 8134 14960 8186
rect 15012 8134 15024 8186
rect 15076 8134 16836 8186
rect 1104 8112 16836 8134
rect 1946 8072 1952 8084
rect 1504 8044 1952 8072
rect 1504 7945 1532 8044
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 4062 8072 4068 8084
rect 2372 8044 4068 8072
rect 2372 8032 2378 8044
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 6178 8072 6184 8084
rect 4172 8044 6184 8072
rect 4172 8004 4200 8044
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 7834 8032 7840 8084
rect 7892 8072 7898 8084
rect 10778 8072 10784 8084
rect 7892 8044 9996 8072
rect 7892 8032 7898 8044
rect 2792 7976 4200 8004
rect 1489 7939 1547 7945
rect 1489 7905 1501 7939
rect 1535 7905 1547 7939
rect 1489 7899 1547 7905
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7936 1823 7939
rect 2792 7936 2820 7976
rect 4430 7964 4436 8016
rect 4488 8004 4494 8016
rect 6733 8007 6791 8013
rect 6733 8004 6745 8007
rect 4488 7976 6745 8004
rect 4488 7964 4494 7976
rect 6733 7973 6745 7976
rect 6779 8004 6791 8007
rect 9968 8004 9996 8044
rect 10152 8044 10784 8072
rect 10152 8004 10180 8044
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 11974 8032 11980 8084
rect 12032 8072 12038 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 12032 8044 15117 8072
rect 12032 8032 12038 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 13354 8004 13360 8016
rect 6779 7976 9904 8004
rect 9968 7976 10180 8004
rect 10244 7976 13360 8004
rect 6779 7973 6791 7976
rect 6733 7967 6791 7973
rect 9398 7936 9404 7948
rect 1811 7908 2820 7936
rect 2884 7908 9168 7936
rect 1811 7905 1823 7908
rect 1765 7899 1823 7905
rect 2884 7854 2912 7908
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 5074 7868 5080 7880
rect 4111 7840 5080 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 3804 7800 3832 7831
rect 5074 7828 5080 7840
rect 5132 7828 5138 7880
rect 7466 7868 7472 7880
rect 7427 7840 7472 7868
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 7558 7828 7564 7880
rect 7616 7868 7622 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7616 7840 7665 7868
rect 7616 7828 7622 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8018 7868 8024 7880
rect 7975 7840 8024 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 4798 7800 4804 7812
rect 3804 7772 4804 7800
rect 4798 7760 4804 7772
rect 4856 7760 4862 7812
rect 5261 7803 5319 7809
rect 5261 7769 5273 7803
rect 5307 7800 5319 7803
rect 8386 7800 8392 7812
rect 5307 7772 8392 7800
rect 5307 7769 5319 7772
rect 5261 7763 5319 7769
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 9140 7800 9168 7908
rect 9232 7908 9404 7936
rect 9232 7880 9260 7908
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 9585 7939 9643 7945
rect 9585 7905 9597 7939
rect 9631 7936 9643 7939
rect 9766 7936 9772 7948
rect 9631 7908 9772 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 9876 7936 9904 7976
rect 10244 7936 10272 7976
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 13538 7964 13544 8016
rect 13596 8004 13602 8016
rect 13596 7976 14320 8004
rect 13596 7964 13602 7976
rect 9876 7908 10272 7936
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 12342 7936 12348 7948
rect 11388 7908 12348 7936
rect 11388 7896 11394 7908
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 12444 7908 13860 7936
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9306 7828 9312 7880
rect 9364 7868 9370 7880
rect 12444 7868 12472 7908
rect 9364 7840 12472 7868
rect 12621 7871 12679 7877
rect 9364 7828 9370 7840
rect 12621 7837 12633 7871
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7868 12955 7871
rect 13446 7868 13452 7880
rect 12943 7840 13452 7868
rect 12943 7837 12955 7840
rect 12897 7831 12955 7837
rect 10410 7800 10416 7812
rect 9140 7772 9987 7800
rect 10371 7772 10416 7800
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 3237 7735 3295 7741
rect 3237 7732 3249 7735
rect 2556 7704 3249 7732
rect 2556 7692 2562 7704
rect 3237 7701 3249 7704
rect 3283 7732 3295 7735
rect 3326 7732 3332 7744
rect 3283 7704 3332 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 3326 7692 3332 7704
rect 3384 7692 3390 7744
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 4614 7732 4620 7744
rect 4212 7704 4620 7732
rect 4212 7692 4218 7704
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 7282 7732 7288 7744
rect 5408 7704 7288 7732
rect 5408 7692 5414 7704
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7837 7735 7895 7741
rect 7837 7701 7849 7735
rect 7883 7732 7895 7735
rect 7926 7732 7932 7744
rect 7883 7704 7932 7732
rect 7883 7701 7895 7704
rect 7837 7695 7895 7701
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8720 7704 8953 7732
rect 8720 7692 8726 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 8941 7695 8999 7701
rect 9030 7692 9036 7744
rect 9088 7732 9094 7744
rect 9309 7735 9367 7741
rect 9309 7732 9321 7735
rect 9088 7704 9321 7732
rect 9088 7692 9094 7704
rect 9309 7701 9321 7704
rect 9355 7701 9367 7735
rect 9309 7695 9367 7701
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 9858 7732 9864 7744
rect 9447 7704 9864 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 9959 7732 9987 7772
rect 10410 7760 10416 7772
rect 10468 7760 10474 7812
rect 10594 7760 10600 7812
rect 10652 7800 10658 7812
rect 10778 7800 10784 7812
rect 10652 7772 10784 7800
rect 10652 7760 10658 7772
rect 10778 7760 10784 7772
rect 10836 7800 10842 7812
rect 12636 7800 12664 7831
rect 13446 7828 13452 7840
rect 13504 7828 13510 7880
rect 13722 7800 13728 7812
rect 10836 7772 13728 7800
rect 10836 7760 10842 7772
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 13832 7800 13860 7908
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 13964 7908 14197 7936
rect 13964 7896 13970 7908
rect 14185 7905 14197 7908
rect 14231 7905 14243 7939
rect 14185 7899 14243 7905
rect 14292 7877 14320 7976
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 14792 7840 15301 7868
rect 14792 7828 14798 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 15378 7828 15384 7880
rect 15436 7868 15442 7880
rect 15473 7871 15531 7877
rect 15473 7868 15485 7871
rect 15436 7840 15485 7868
rect 15436 7828 15442 7840
rect 15473 7837 15485 7840
rect 15519 7837 15531 7871
rect 15473 7831 15531 7837
rect 15565 7871 15623 7877
rect 15565 7837 15577 7871
rect 15611 7868 15623 7871
rect 16206 7868 16212 7880
rect 15611 7840 16212 7868
rect 15611 7837 15623 7840
rect 15565 7831 15623 7837
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 16666 7800 16672 7812
rect 13832 7772 16672 7800
rect 16666 7760 16672 7772
rect 16724 7760 16730 7812
rect 11330 7732 11336 7744
rect 9959 7704 11336 7732
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 11514 7692 11520 7744
rect 11572 7732 11578 7744
rect 11701 7735 11759 7741
rect 11701 7732 11713 7735
rect 11572 7704 11713 7732
rect 11572 7692 11578 7704
rect 11701 7701 11713 7704
rect 11747 7701 11759 7735
rect 11701 7695 11759 7701
rect 11974 7692 11980 7744
rect 12032 7732 12038 7744
rect 13906 7732 13912 7744
rect 12032 7704 13912 7732
rect 12032 7692 12038 7704
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 14642 7732 14648 7744
rect 14603 7704 14648 7732
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 16390 7732 16396 7744
rect 14884 7704 16396 7732
rect 14884 7692 14890 7704
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 1104 7642 16836 7664
rect 1104 7590 4898 7642
rect 4950 7590 4962 7642
rect 5014 7590 5026 7642
rect 5078 7590 5090 7642
rect 5142 7590 5154 7642
rect 5206 7590 8846 7642
rect 8898 7590 8910 7642
rect 8962 7590 8974 7642
rect 9026 7590 9038 7642
rect 9090 7590 9102 7642
rect 9154 7590 12794 7642
rect 12846 7590 12858 7642
rect 12910 7590 12922 7642
rect 12974 7590 12986 7642
rect 13038 7590 13050 7642
rect 13102 7590 16836 7642
rect 1104 7568 16836 7590
rect 1946 7488 1952 7540
rect 2004 7488 2010 7540
rect 9490 7528 9496 7540
rect 4080 7500 9496 7528
rect 1964 7460 1992 7488
rect 4080 7469 4108 7500
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 11422 7528 11428 7540
rect 10152 7500 11428 7528
rect 1872 7432 1992 7460
rect 4065 7463 4123 7469
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 1872 7401 1900 7432
rect 4065 7429 4077 7463
rect 4111 7429 4123 7463
rect 4065 7423 4123 7429
rect 5813 7463 5871 7469
rect 5813 7429 5825 7463
rect 5859 7460 5871 7463
rect 7374 7460 7380 7472
rect 5859 7432 7380 7460
rect 5859 7429 5871 7432
rect 5813 7423 5871 7429
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 7834 7460 7840 7472
rect 7795 7432 7840 7460
rect 7834 7420 7840 7432
rect 7892 7420 7898 7472
rect 7926 7420 7932 7472
rect 7984 7460 7990 7472
rect 10152 7460 10180 7500
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 12066 7488 12072 7540
rect 12124 7528 12130 7540
rect 12894 7528 12900 7540
rect 12124 7500 12900 7528
rect 12124 7488 12130 7500
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 13906 7528 13912 7540
rect 13286 7500 13912 7528
rect 11974 7460 11980 7472
rect 7984 7432 10180 7460
rect 10796 7432 11980 7460
rect 7984 7420 7990 7432
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1544 7364 1869 7392
rect 1544 7352 1550 7364
rect 1857 7361 1869 7364
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7324 2191 7327
rect 2682 7324 2688 7336
rect 2179 7296 2688 7324
rect 2179 7293 2191 7296
rect 2133 7287 2191 7293
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 3252 7256 3280 7378
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 7006 7392 7012 7404
rect 6052 7364 7012 7392
rect 6052 7352 6058 7364
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7101 7395 7159 7401
rect 7101 7361 7113 7395
rect 7147 7392 7159 7395
rect 7742 7392 7748 7404
rect 7147 7364 7748 7392
rect 7147 7361 7159 7364
rect 7101 7355 7159 7361
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 10594 7392 10600 7404
rect 10555 7364 10600 7392
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 6270 7324 6276 7336
rect 5684 7296 6276 7324
rect 5684 7284 5690 7296
rect 6270 7284 6276 7296
rect 6328 7324 6334 7336
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 6328 7296 7205 7324
rect 6328 7284 6334 7296
rect 7193 7293 7205 7296
rect 7239 7293 7251 7327
rect 7193 7287 7251 7293
rect 7282 7284 7288 7336
rect 7340 7324 7346 7336
rect 10796 7333 10824 7432
rect 11974 7420 11980 7432
rect 12032 7420 12038 7472
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 12621 7463 12679 7469
rect 12621 7460 12633 7463
rect 12584 7432 12633 7460
rect 12584 7420 12590 7432
rect 12621 7429 12633 7432
rect 12667 7429 12679 7463
rect 13286 7460 13314 7500
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 15378 7488 15384 7540
rect 15436 7528 15442 7540
rect 16942 7528 16948 7540
rect 15436 7500 16948 7528
rect 15436 7488 15442 7500
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 12621 7423 12679 7429
rect 12912 7432 13314 7460
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7361 10931 7395
rect 10873 7355 10931 7361
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 11882 7392 11888 7404
rect 11839 7364 11888 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 7340 7296 10793 7324
rect 7340 7284 7346 7296
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 10888 7324 10916 7355
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7392 12127 7395
rect 12636 7392 12756 7393
rect 12912 7392 12940 7432
rect 13354 7420 13360 7472
rect 13412 7460 13418 7472
rect 14734 7460 14740 7472
rect 13412 7432 14740 7460
rect 13412 7420 13418 7432
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 15010 7420 15016 7472
rect 15068 7460 15074 7472
rect 15068 7432 15608 7460
rect 15068 7420 15074 7432
rect 12115 7372 12572 7392
rect 12636 7372 12940 7392
rect 12115 7365 12940 7372
rect 12115 7364 12664 7365
rect 12728 7364 12940 7365
rect 12115 7361 12127 7364
rect 12069 7355 12127 7361
rect 12544 7344 12664 7364
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 14826 7392 14832 7404
rect 13044 7364 14832 7392
rect 13044 7352 13050 7364
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7361 15347 7395
rect 15289 7355 15347 7361
rect 11238 7324 11244 7336
rect 10888 7296 11244 7324
rect 10781 7287 10839 7293
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7324 11759 7327
rect 11974 7324 11980 7336
rect 11747 7296 11980 7324
rect 11747 7293 11759 7296
rect 11701 7287 11759 7293
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7324 12219 7327
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 12207 7296 12480 7324
rect 12207 7293 12219 7296
rect 12161 7287 12219 7293
rect 7926 7256 7932 7268
rect 3252 7228 7932 7256
rect 7926 7216 7932 7228
rect 7984 7216 7990 7268
rect 8938 7216 8944 7268
rect 8996 7256 9002 7268
rect 9766 7256 9772 7268
rect 8996 7228 9772 7256
rect 8996 7216 9002 7228
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 10686 7256 10692 7268
rect 10647 7228 10692 7256
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 11517 7259 11575 7265
rect 11517 7225 11529 7259
rect 11563 7256 11575 7259
rect 11606 7256 11612 7268
rect 11563 7228 11612 7256
rect 11563 7225 11575 7228
rect 11517 7219 11575 7225
rect 11606 7216 11612 7228
rect 11664 7216 11670 7268
rect 12452 7256 12480 7296
rect 12728 7296 15117 7324
rect 12728 7256 12756 7296
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15304 7324 15332 7355
rect 15378 7352 15384 7404
rect 15436 7392 15442 7404
rect 15580 7401 15608 7432
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15436 7364 15485 7392
rect 15436 7352 15442 7364
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7361 15623 7395
rect 15565 7355 15623 7361
rect 15304 7296 15608 7324
rect 15105 7287 15163 7293
rect 15580 7268 15608 7296
rect 12452 7228 12756 7256
rect 12802 7216 12808 7268
rect 12860 7256 12866 7268
rect 12860 7228 15516 7256
rect 12860 7216 12866 7228
rect 3605 7191 3663 7197
rect 3605 7157 3617 7191
rect 3651 7188 3663 7191
rect 3694 7188 3700 7200
rect 3651 7160 3700 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 3694 7148 3700 7160
rect 3752 7148 3758 7200
rect 4062 7148 4068 7200
rect 4120 7188 4126 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 4120 7160 6653 7188
rect 4120 7148 4126 7160
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 6641 7151 6699 7157
rect 7466 7148 7472 7200
rect 7524 7188 7530 7200
rect 8386 7188 8392 7200
rect 7524 7160 8392 7188
rect 7524 7148 7530 7160
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 8628 7160 9137 7188
rect 8628 7148 8634 7160
rect 9125 7157 9137 7160
rect 9171 7188 9183 7191
rect 9582 7188 9588 7200
rect 9171 7160 9588 7188
rect 9171 7157 9183 7160
rect 9125 7151 9183 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 10413 7191 10471 7197
rect 10413 7157 10425 7191
rect 10459 7188 10471 7191
rect 12710 7188 12716 7200
rect 10459 7160 12716 7188
rect 10459 7157 10471 7160
rect 10413 7151 10471 7157
rect 12710 7148 12716 7160
rect 12768 7148 12774 7200
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13909 7191 13967 7197
rect 13909 7188 13921 7191
rect 13228 7160 13921 7188
rect 13228 7148 13234 7160
rect 13909 7157 13921 7160
rect 13955 7157 13967 7191
rect 15488 7188 15516 7228
rect 15562 7216 15568 7268
rect 15620 7256 15626 7268
rect 15746 7256 15752 7268
rect 15620 7228 15752 7256
rect 15620 7216 15626 7228
rect 15746 7216 15752 7228
rect 15804 7216 15810 7268
rect 16206 7188 16212 7200
rect 15488 7160 16212 7188
rect 13909 7151 13967 7157
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 1104 7098 16836 7120
rect 1104 7046 2924 7098
rect 2976 7046 2988 7098
rect 3040 7046 3052 7098
rect 3104 7046 3116 7098
rect 3168 7046 3180 7098
rect 3232 7046 6872 7098
rect 6924 7046 6936 7098
rect 6988 7046 7000 7098
rect 7052 7046 7064 7098
rect 7116 7046 7128 7098
rect 7180 7046 10820 7098
rect 10872 7046 10884 7098
rect 10936 7046 10948 7098
rect 11000 7046 11012 7098
rect 11064 7046 11076 7098
rect 11128 7046 14768 7098
rect 14820 7046 14832 7098
rect 14884 7046 14896 7098
rect 14948 7046 14960 7098
rect 15012 7046 15024 7098
rect 15076 7046 16836 7098
rect 1104 7024 16836 7046
rect 1752 6987 1810 6993
rect 1752 6953 1764 6987
rect 1798 6984 1810 6987
rect 2222 6984 2228 6996
rect 1798 6956 2228 6984
rect 1798 6953 1810 6956
rect 1752 6947 1810 6953
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 4080 6956 4476 6984
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 4080 6848 4108 6956
rect 4338 6848 4344 6860
rect 1820 6820 4108 6848
rect 4172 6820 4344 6848
rect 1820 6808 1826 6820
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6780 4031 6783
rect 4172 6780 4200 6820
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 4448 6848 4476 6956
rect 7466 6944 7472 6996
rect 7524 6984 7530 6996
rect 7524 6956 8708 6984
rect 7524 6944 7530 6956
rect 5166 6876 5172 6928
rect 5224 6916 5230 6928
rect 7558 6916 7564 6928
rect 5224 6888 7564 6916
rect 5224 6876 5230 6888
rect 7558 6876 7564 6888
rect 7616 6876 7622 6928
rect 8680 6916 8708 6956
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 9582 6984 9588 6996
rect 8812 6956 9588 6984
rect 8812 6944 8818 6956
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 11057 6987 11115 6993
rect 9681 6956 10732 6984
rect 9125 6919 9183 6925
rect 9125 6916 9137 6919
rect 7659 6888 8524 6916
rect 8680 6888 9137 6916
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 4448 6820 6837 6848
rect 6825 6817 6837 6820
rect 6871 6817 6883 6851
rect 6825 6811 6883 6817
rect 4019 6752 4200 6780
rect 4249 6783 4307 6789
rect 4019 6749 4031 6752
rect 3973 6743 4031 6749
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 5166 6780 5172 6792
rect 4295 6752 5172 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6780 5319 6783
rect 5442 6780 5448 6792
rect 5307 6752 5448 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 7659 6780 7687 6888
rect 7834 6808 7840 6860
rect 7892 6848 7898 6860
rect 7892 6820 8248 6848
rect 7892 6808 7898 6820
rect 8018 6780 8024 6792
rect 5552 6752 7687 6780
rect 7979 6752 8024 6780
rect 4798 6712 4804 6724
rect 2990 6684 4804 6712
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 4062 6644 4068 6656
rect 3283 6616 4068 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 4614 6604 4620 6656
rect 4672 6644 4678 6656
rect 5552 6644 5580 6752
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8220 6789 8248 6820
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 6454 6672 6460 6724
rect 6512 6712 6518 6724
rect 8389 6715 8447 6721
rect 8389 6712 8401 6715
rect 6512 6684 8401 6712
rect 6512 6672 6518 6684
rect 8389 6681 8401 6684
rect 8435 6681 8447 6715
rect 8496 6712 8524 6888
rect 9125 6885 9137 6888
rect 9171 6885 9183 6919
rect 9681 6916 9709 6956
rect 9125 6879 9183 6885
rect 9416 6888 9709 6916
rect 9416 6860 9444 6888
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9217 6851 9275 6857
rect 9217 6848 9229 6851
rect 8904 6820 9229 6848
rect 8904 6808 8910 6820
rect 9217 6817 9229 6820
rect 9263 6817 9275 6851
rect 9217 6811 9275 6817
rect 9398 6808 9404 6860
rect 9456 6808 9462 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9499 6820 9689 6848
rect 8938 6780 8944 6792
rect 8899 6752 8944 6780
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9033 6783 9091 6789
rect 9033 6749 9045 6783
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9048 6712 9076 6743
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9499 6780 9527 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 10704 6848 10732 6956
rect 11057 6953 11069 6987
rect 11103 6984 11115 6987
rect 11422 6984 11428 6996
rect 11103 6956 11428 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 11422 6944 11428 6956
rect 11480 6984 11486 6996
rect 13262 6984 13268 6996
rect 11480 6956 13268 6984
rect 11480 6944 11486 6956
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 14734 6944 14740 6996
rect 14792 6984 14798 6996
rect 16298 6984 16304 6996
rect 14792 6956 16304 6984
rect 14792 6944 14798 6956
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 12618 6876 12624 6928
rect 12676 6916 12682 6928
rect 12897 6919 12955 6925
rect 12897 6916 12909 6919
rect 12676 6888 12909 6916
rect 12676 6876 12682 6888
rect 12897 6885 12909 6888
rect 12943 6885 12955 6919
rect 12897 6879 12955 6885
rect 13188 6888 14412 6916
rect 10704 6820 11652 6848
rect 9677 6811 9735 6817
rect 11624 6792 11652 6820
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 13188 6848 13216 6888
rect 14384 6848 14412 6888
rect 15194 6876 15200 6928
rect 15252 6876 15258 6928
rect 15289 6919 15347 6925
rect 15289 6885 15301 6919
rect 15335 6916 15347 6919
rect 16666 6916 16672 6928
rect 15335 6888 16672 6916
rect 15335 6885 15347 6888
rect 15289 6879 15347 6885
rect 16666 6876 16672 6888
rect 16724 6876 16730 6928
rect 15212 6848 15240 6876
rect 12584 6820 13216 6848
rect 13280 6820 14320 6848
rect 14384 6820 15056 6848
rect 15212 6820 16160 6848
rect 12584 6808 12590 6820
rect 9364 6752 9527 6780
rect 9944 6783 10002 6789
rect 9364 6740 9370 6752
rect 9944 6749 9956 6783
rect 9990 6780 10002 6783
rect 10778 6782 10784 6792
rect 10704 6780 10784 6782
rect 9990 6754 10784 6780
rect 9990 6752 10732 6754
rect 9990 6749 10002 6752
rect 9944 6743 10002 6749
rect 10778 6740 10784 6754
rect 10836 6740 10842 6792
rect 10870 6740 10876 6792
rect 10928 6780 10934 6792
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 10928 6752 11529 6780
rect 10928 6740 10934 6752
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 11606 6740 11612 6792
rect 11664 6740 11670 6792
rect 11784 6783 11842 6789
rect 11784 6749 11796 6783
rect 11830 6780 11842 6783
rect 12250 6780 12256 6792
rect 11830 6752 12256 6780
rect 11830 6749 11842 6752
rect 11784 6743 11842 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 12894 6740 12900 6792
rect 12952 6780 12958 6792
rect 13280 6780 13308 6820
rect 12952 6752 13308 6780
rect 12952 6740 12958 6752
rect 13354 6740 13360 6792
rect 13412 6780 13418 6792
rect 14093 6783 14151 6789
rect 13412 6752 13457 6780
rect 13412 6740 13418 6752
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 14182 6780 14188 6792
rect 14139 6752 14188 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 14182 6740 14188 6752
rect 14240 6740 14246 6792
rect 14292 6789 14320 6820
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 14734 6780 14740 6792
rect 14599 6752 14740 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 15028 6789 15056 6820
rect 15194 6789 15200 6792
rect 15013 6783 15071 6789
rect 15013 6749 15025 6783
rect 15059 6749 15071 6783
rect 15013 6743 15071 6749
rect 15151 6783 15200 6789
rect 15151 6749 15163 6783
rect 15197 6749 15200 6783
rect 15151 6743 15200 6749
rect 15194 6740 15200 6743
rect 15252 6740 15258 6792
rect 15470 6780 15476 6792
rect 15431 6752 15476 6780
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 16132 6789 16160 6820
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 8496 6684 9076 6712
rect 8389 6675 8447 6681
rect 9122 6672 9128 6724
rect 9180 6712 9186 6724
rect 11422 6712 11428 6724
rect 9180 6684 11428 6712
rect 9180 6672 9186 6684
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 15381 6715 15439 6721
rect 15381 6712 15393 6715
rect 11532 6684 15393 6712
rect 4672 6616 5580 6644
rect 4672 6604 4678 6616
rect 6730 6604 6736 6656
rect 6788 6644 6794 6656
rect 9582 6644 9588 6656
rect 6788 6616 9588 6644
rect 6788 6604 6794 6616
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 10042 6604 10048 6656
rect 10100 6644 10106 6656
rect 10686 6644 10692 6656
rect 10100 6616 10692 6644
rect 10100 6604 10106 6616
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 11532 6644 11560 6684
rect 15381 6681 15393 6684
rect 15427 6681 15439 6715
rect 15381 6675 15439 6681
rect 10836 6616 11560 6644
rect 10836 6604 10842 6616
rect 11974 6604 11980 6656
rect 12032 6644 12038 6656
rect 12526 6644 12532 6656
rect 12032 6616 12532 6644
rect 12032 6604 12038 6616
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 13446 6644 13452 6656
rect 13407 6616 13452 6644
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 13872 6616 14473 6644
rect 13872 6604 13878 6616
rect 14461 6613 14473 6616
rect 14507 6613 14519 6647
rect 14461 6607 14519 6613
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 15933 6647 15991 6653
rect 15933 6644 15945 6647
rect 15620 6616 15945 6644
rect 15620 6604 15626 6616
rect 15933 6613 15945 6616
rect 15979 6613 15991 6647
rect 15933 6607 15991 6613
rect 1104 6554 16836 6576
rect 1104 6502 4898 6554
rect 4950 6502 4962 6554
rect 5014 6502 5026 6554
rect 5078 6502 5090 6554
rect 5142 6502 5154 6554
rect 5206 6502 8846 6554
rect 8898 6502 8910 6554
rect 8962 6502 8974 6554
rect 9026 6502 9038 6554
rect 9090 6502 9102 6554
rect 9154 6502 12794 6554
rect 12846 6502 12858 6554
rect 12910 6502 12922 6554
rect 12974 6502 12986 6554
rect 13038 6502 13050 6554
rect 13102 6502 16836 6554
rect 1104 6480 16836 6502
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 5537 6443 5595 6449
rect 5537 6440 5549 6443
rect 2832 6412 5549 6440
rect 2832 6400 2838 6412
rect 5537 6409 5549 6412
rect 5583 6409 5595 6443
rect 5537 6403 5595 6409
rect 6917 6443 6975 6449
rect 6917 6409 6929 6443
rect 6963 6440 6975 6443
rect 7650 6440 7656 6452
rect 6963 6412 7656 6440
rect 6963 6409 6975 6412
rect 6917 6403 6975 6409
rect 7650 6400 7656 6412
rect 7708 6400 7714 6452
rect 8754 6440 8760 6452
rect 8715 6412 8760 6440
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 10410 6440 10416 6452
rect 9159 6412 10416 6440
rect 4338 6372 4344 6384
rect 3082 6344 4344 6372
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 8202 6372 8208 6384
rect 5290 6344 8208 6372
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1544 6276 1593 6304
rect 1544 6264 1550 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 5902 6264 5908 6316
rect 5960 6304 5966 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5960 6276 6377 6304
rect 5960 6264 5966 6276
rect 6365 6273 6377 6276
rect 6411 6304 6423 6307
rect 6454 6304 6460 6316
rect 6411 6276 6460 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6304 6791 6307
rect 7098 6304 7104 6316
rect 6779 6276 7104 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 3694 6236 3700 6248
rect 1903 6208 3700 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 3694 6196 3700 6208
rect 3752 6196 3758 6248
rect 3789 6239 3847 6245
rect 3789 6205 3801 6239
rect 3835 6236 3847 6239
rect 4065 6239 4123 6245
rect 3835 6208 3924 6236
rect 3835 6205 3847 6208
rect 3789 6199 3847 6205
rect 3896 6168 3924 6208
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 5350 6236 5356 6248
rect 4111 6208 5356 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 5810 6236 5816 6248
rect 5592 6208 5816 6236
rect 5592 6196 5598 6208
rect 5810 6196 5816 6208
rect 5868 6236 5874 6248
rect 6564 6236 6592 6267
rect 5868 6208 6592 6236
rect 5868 6196 5874 6208
rect 3252 6140 3924 6168
rect 6656 6168 6684 6267
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7374 6304 7380 6316
rect 7248 6276 7380 6304
rect 7248 6264 7254 6276
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 7644 6307 7702 6313
rect 7644 6273 7656 6307
rect 7690 6304 7702 6307
rect 9159 6304 9187 6412
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 14737 6443 14795 6449
rect 14737 6440 14749 6443
rect 13136 6412 14749 6440
rect 13136 6400 13142 6412
rect 14737 6409 14749 6412
rect 14783 6409 14795 6443
rect 14737 6403 14795 6409
rect 11514 6372 11520 6384
rect 9232 6344 11520 6372
rect 9232 6313 9260 6344
rect 11514 6332 11520 6344
rect 11572 6332 11578 6384
rect 11974 6332 11980 6384
rect 12032 6372 12038 6384
rect 14277 6375 14335 6381
rect 12032 6344 13860 6372
rect 12032 6332 12038 6344
rect 7690 6276 9187 6304
rect 9217 6307 9275 6313
rect 7690 6273 7702 6276
rect 7644 6267 7702 6273
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 9484 6307 9542 6313
rect 9484 6273 9496 6307
rect 9530 6304 9542 6307
rect 11146 6304 11152 6316
rect 9530 6276 11152 6304
rect 9530 6273 9542 6276
rect 9484 6267 9542 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11773 6307 11831 6313
rect 11773 6304 11785 6307
rect 11256 6276 11785 6304
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 9324 6236 9352 6264
rect 8996 6208 9352 6236
rect 8996 6196 9002 6208
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 11256 6236 11284 6276
rect 11773 6273 11785 6276
rect 11819 6273 11831 6307
rect 11773 6267 11831 6273
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 13832 6313 13860 6344
rect 14277 6341 14289 6375
rect 14323 6372 14335 6375
rect 14642 6372 14648 6384
rect 14323 6344 14648 6372
rect 14323 6341 14335 6344
rect 14277 6335 14335 6341
rect 14642 6332 14648 6344
rect 14700 6332 14706 6384
rect 17494 6372 17500 6384
rect 15212 6344 17500 6372
rect 13541 6307 13599 6313
rect 13541 6304 13553 6307
rect 13412 6276 13553 6304
rect 13412 6264 13418 6276
rect 13541 6273 13553 6276
rect 13587 6273 13599 6307
rect 13541 6267 13599 6273
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 11514 6236 11520 6248
rect 10376 6208 11284 6236
rect 11475 6208 11520 6236
rect 10376 6196 10382 6208
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 7374 6168 7380 6180
rect 6656 6140 7380 6168
rect 1486 6060 1492 6112
rect 1544 6100 1550 6112
rect 3252 6100 3280 6140
rect 1544 6072 3280 6100
rect 1544 6060 1550 6072
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3896 6100 3924 6140
rect 7374 6128 7380 6140
rect 7432 6128 7438 6180
rect 8312 6140 8892 6168
rect 5350 6100 5356 6112
rect 3384 6072 3429 6100
rect 3896 6072 5356 6100
rect 3384 6060 3390 6072
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 6546 6060 6552 6112
rect 6604 6100 6610 6112
rect 8312 6100 8340 6140
rect 6604 6072 8340 6100
rect 8864 6100 8892 6140
rect 10152 6140 10732 6168
rect 10152 6100 10180 6140
rect 8864 6072 10180 6100
rect 6604 6060 6610 6072
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 10376 6072 10609 6100
rect 10376 6060 10382 6072
rect 10597 6069 10609 6072
rect 10643 6069 10655 6103
rect 10704 6100 10732 6140
rect 12710 6128 12716 6180
rect 12768 6168 12774 6180
rect 13357 6171 13415 6177
rect 13357 6168 13369 6171
rect 12768 6140 13369 6168
rect 12768 6128 12774 6140
rect 13357 6137 13369 6140
rect 13403 6137 13415 6171
rect 13357 6131 13415 6137
rect 12158 6100 12164 6112
rect 10704 6072 12164 6100
rect 10597 6063 10655 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12526 6060 12532 6112
rect 12584 6100 12590 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 12584 6072 12909 6100
rect 12584 6060 12590 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 12897 6063 12955 6069
rect 13262 6060 13268 6112
rect 13320 6100 13326 6112
rect 13538 6100 13544 6112
rect 13320 6072 13544 6100
rect 13320 6060 13326 6072
rect 13538 6060 13544 6072
rect 13596 6100 13602 6112
rect 13740 6100 13768 6267
rect 14550 6264 14556 6316
rect 14608 6264 14614 6316
rect 15212 6313 15240 6344
rect 17494 6332 17500 6344
rect 17552 6332 17558 6384
rect 15197 6307 15255 6313
rect 15197 6273 15209 6307
rect 15243 6273 15255 6307
rect 15197 6267 15255 6273
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6304 15439 6307
rect 17126 6304 17132 6316
rect 15427 6276 17132 6304
rect 15427 6273 15439 6276
rect 15381 6267 15439 6273
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 14568 6236 14596 6264
rect 14568 6208 15148 6236
rect 14090 6128 14096 6180
rect 14148 6168 14154 6180
rect 14553 6171 14611 6177
rect 14553 6168 14565 6171
rect 14148 6140 14565 6168
rect 14148 6128 14154 6140
rect 14553 6137 14565 6140
rect 14599 6137 14611 6171
rect 14553 6131 14611 6137
rect 13596 6072 13768 6100
rect 15120 6100 15148 6208
rect 15197 6103 15255 6109
rect 15197 6100 15209 6103
rect 15120 6072 15209 6100
rect 13596 6060 13602 6072
rect 15197 6069 15209 6072
rect 15243 6069 15255 6103
rect 15562 6100 15568 6112
rect 15523 6072 15568 6100
rect 15197 6063 15255 6069
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 1104 6010 16836 6032
rect 1104 5958 2924 6010
rect 2976 5958 2988 6010
rect 3040 5958 3052 6010
rect 3104 5958 3116 6010
rect 3168 5958 3180 6010
rect 3232 5958 6872 6010
rect 6924 5958 6936 6010
rect 6988 5958 7000 6010
rect 7052 5958 7064 6010
rect 7116 5958 7128 6010
rect 7180 5958 10820 6010
rect 10872 5958 10884 6010
rect 10936 5958 10948 6010
rect 11000 5958 11012 6010
rect 11064 5958 11076 6010
rect 11128 5958 14768 6010
rect 14820 5958 14832 6010
rect 14884 5958 14896 6010
rect 14948 5958 14960 6010
rect 15012 5958 15024 6010
rect 15076 5958 16836 6010
rect 1104 5936 16836 5958
rect 6546 5896 6552 5908
rect 3252 5868 6552 5896
rect 1486 5760 1492 5772
rect 1447 5732 1492 5760
rect 1486 5720 1492 5732
rect 1544 5720 1550 5772
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 3252 5760 3280 5868
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 6730 5896 6736 5908
rect 6691 5868 6736 5896
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7834 5896 7840 5908
rect 7432 5868 7840 5896
rect 7432 5856 7438 5868
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 7926 5856 7932 5908
rect 7984 5896 7990 5908
rect 9309 5899 9367 5905
rect 7984 5868 9260 5896
rect 7984 5856 7990 5868
rect 3326 5788 3332 5840
rect 3384 5828 3390 5840
rect 8846 5828 8852 5840
rect 3384 5800 8852 5828
rect 3384 5788 3390 5800
rect 8846 5788 8852 5800
rect 8904 5788 8910 5840
rect 9232 5828 9260 5868
rect 9309 5865 9321 5899
rect 9355 5896 9367 5899
rect 11882 5896 11888 5908
rect 9355 5868 11008 5896
rect 9355 5865 9367 5868
rect 9309 5859 9367 5865
rect 9674 5828 9680 5840
rect 9232 5800 9680 5828
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 9784 5800 10180 5828
rect 3510 5760 3516 5772
rect 1811 5732 3280 5760
rect 3344 5732 3516 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 3344 5704 3372 5732
rect 3510 5720 3516 5732
rect 3568 5760 3574 5772
rect 3973 5763 4031 5769
rect 3973 5760 3985 5763
rect 3568 5732 3985 5760
rect 3568 5720 3574 5732
rect 3973 5729 3985 5732
rect 4019 5729 4031 5763
rect 6638 5760 6644 5772
rect 3973 5723 4031 5729
rect 5276 5732 6644 5760
rect 3326 5652 3332 5704
rect 3384 5652 3390 5704
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 5276 5701 5304 5732
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 8478 5760 8484 5772
rect 8036 5732 8484 5760
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 4120 5664 4261 5692
rect 4120 5652 4126 5664
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5661 5319 5695
rect 5261 5655 5319 5661
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 7926 5692 7932 5704
rect 5592 5664 7932 5692
rect 5592 5652 5598 5664
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 8036 5701 8064 5732
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 9784 5760 9812 5800
rect 9508 5732 9812 5760
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8110 5652 8116 5704
rect 8168 5692 8174 5704
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 8168 5664 8217 5692
rect 8168 5652 8174 5664
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 9214 5692 9220 5704
rect 8343 5664 9220 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9508 5701 9536 5732
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 9766 5652 9772 5704
rect 9824 5701 9830 5704
rect 9824 5695 9873 5701
rect 9824 5661 9827 5695
rect 9861 5661 9873 5695
rect 9824 5655 9873 5661
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 9824 5652 9830 5655
rect 2990 5596 8432 5624
rect 2038 5516 2044 5568
rect 2096 5556 2102 5568
rect 2774 5556 2780 5568
rect 2096 5528 2780 5556
rect 2096 5516 2102 5528
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 3510 5556 3516 5568
rect 3283 5528 3516 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 3510 5516 3516 5528
rect 3568 5516 3574 5568
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 4062 5556 4068 5568
rect 3752 5528 4068 5556
rect 3752 5516 3758 5528
rect 4062 5516 4068 5528
rect 4120 5556 4126 5568
rect 7650 5556 7656 5568
rect 4120 5528 7656 5556
rect 4120 5516 4126 5528
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 7837 5559 7895 5565
rect 7837 5525 7849 5559
rect 7883 5556 7895 5559
rect 8110 5556 8116 5568
rect 7883 5528 8116 5556
rect 7883 5525 7895 5528
rect 7837 5519 7895 5525
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8404 5556 8432 5596
rect 8478 5584 8484 5636
rect 8536 5624 8542 5636
rect 8536 5596 9168 5624
rect 8536 5584 8542 5596
rect 9030 5556 9036 5568
rect 8404 5528 9036 5556
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 9140 5556 9168 5596
rect 9306 5584 9312 5636
rect 9364 5624 9370 5636
rect 9582 5627 9640 5633
rect 9582 5624 9594 5627
rect 9364 5596 9594 5624
rect 9364 5584 9370 5596
rect 9582 5593 9594 5596
rect 9628 5593 9640 5627
rect 9582 5587 9640 5593
rect 9677 5627 9735 5633
rect 9677 5593 9689 5627
rect 9723 5593 9735 5627
rect 9677 5587 9735 5593
rect 9692 5556 9720 5587
rect 9140 5528 9720 5556
rect 9858 5516 9864 5568
rect 9916 5556 9922 5568
rect 9968 5556 9996 5655
rect 10152 5624 10180 5800
rect 10226 5788 10232 5840
rect 10284 5828 10290 5840
rect 10284 5800 10456 5828
rect 10284 5788 10290 5800
rect 10428 5760 10456 5800
rect 10502 5788 10508 5840
rect 10560 5828 10566 5840
rect 10980 5828 11008 5868
rect 11440 5868 11888 5896
rect 11440 5828 11468 5868
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 13446 5896 13452 5908
rect 12400 5868 13452 5896
rect 12400 5856 12406 5868
rect 13446 5856 13452 5868
rect 13504 5896 13510 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13504 5868 14105 5896
rect 13504 5856 13510 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 14458 5896 14464 5908
rect 14419 5868 14464 5896
rect 14093 5859 14151 5865
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 15102 5856 15108 5908
rect 15160 5896 15166 5908
rect 15841 5899 15899 5905
rect 15841 5896 15853 5899
rect 15160 5868 15853 5896
rect 15160 5856 15166 5868
rect 15841 5865 15853 5868
rect 15887 5865 15899 5899
rect 15841 5859 15899 5865
rect 12434 5828 12440 5840
rect 10560 5800 10916 5828
rect 10980 5800 11468 5828
rect 11532 5800 12440 5828
rect 10560 5788 10566 5800
rect 10778 5760 10784 5772
rect 10428 5732 10784 5760
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 10888 5760 10916 5800
rect 11532 5760 11560 5800
rect 12434 5788 12440 5800
rect 12492 5788 12498 5840
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 15378 5828 15384 5840
rect 12584 5800 15384 5828
rect 12584 5788 12590 5800
rect 15378 5788 15384 5800
rect 15436 5788 15442 5840
rect 11882 5760 11888 5772
rect 10888 5732 11560 5760
rect 11788 5732 11888 5760
rect 11788 5702 11816 5732
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 12618 5720 12624 5772
rect 12676 5760 12682 5772
rect 12989 5763 13047 5769
rect 12989 5760 13001 5763
rect 12676 5732 13001 5760
rect 12676 5720 12682 5732
rect 12989 5729 13001 5732
rect 13035 5729 13047 5763
rect 12989 5723 13047 5729
rect 13078 5720 13084 5772
rect 13136 5760 13142 5772
rect 13538 5760 13544 5772
rect 13136 5732 13544 5760
rect 13136 5720 13142 5732
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 14185 5763 14243 5769
rect 14185 5760 14197 5763
rect 13780 5732 14197 5760
rect 13780 5720 13786 5732
rect 14185 5729 14197 5732
rect 14231 5729 14243 5763
rect 14185 5723 14243 5729
rect 14550 5720 14556 5772
rect 14608 5760 14614 5772
rect 14608 5732 15976 5760
rect 14608 5720 14614 5732
rect 10246 5695 10304 5701
rect 10246 5661 10258 5695
rect 10292 5692 10304 5695
rect 11256 5692 11816 5702
rect 14090 5692 14096 5704
rect 10292 5674 11816 5692
rect 10292 5664 11284 5674
rect 14051 5664 14096 5692
rect 10292 5661 10304 5664
rect 10246 5655 10304 5661
rect 14090 5652 14096 5664
rect 14148 5692 14154 5704
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 14148 5664 15301 5692
rect 14148 5652 14154 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 15838 5692 15844 5704
rect 15799 5664 15844 5692
rect 15289 5655 15347 5661
rect 11606 5624 11612 5636
rect 10152 5596 11612 5624
rect 11606 5584 11612 5596
rect 11664 5584 11670 5636
rect 12621 5627 12679 5633
rect 12621 5624 12633 5627
rect 12268 5596 12633 5624
rect 9916 5528 9996 5556
rect 9916 5516 9922 5528
rect 11422 5516 11428 5568
rect 11480 5556 11486 5568
rect 11517 5559 11575 5565
rect 11517 5556 11529 5559
rect 11480 5528 11529 5556
rect 11480 5516 11486 5528
rect 11517 5525 11529 5528
rect 11563 5525 11575 5559
rect 11517 5519 11575 5525
rect 12066 5516 12072 5568
rect 12124 5556 12130 5568
rect 12268 5565 12296 5596
rect 12621 5593 12633 5596
rect 12667 5593 12679 5627
rect 12802 5624 12808 5636
rect 12763 5596 12808 5624
rect 12621 5587 12679 5593
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 14921 5627 14979 5633
rect 14921 5624 14933 5627
rect 12912 5596 14933 5624
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 12124 5528 12265 5556
rect 12124 5516 12130 5528
rect 12253 5525 12265 5528
rect 12299 5525 12311 5559
rect 12253 5519 12311 5525
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 12912 5556 12940 5596
rect 14921 5593 14933 5596
rect 14967 5593 14979 5627
rect 14921 5587 14979 5593
rect 15105 5627 15163 5633
rect 15105 5593 15117 5627
rect 15151 5593 15163 5627
rect 15304 5624 15332 5655
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 15948 5701 15976 5732
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 16022 5624 16028 5636
rect 15304 5596 16028 5624
rect 15105 5587 15163 5593
rect 12492 5528 12940 5556
rect 12492 5516 12498 5528
rect 13354 5516 13360 5568
rect 13412 5556 13418 5568
rect 15120 5556 15148 5587
rect 16022 5584 16028 5596
rect 16080 5584 16086 5636
rect 13412 5528 15148 5556
rect 13412 5516 13418 5528
rect 1104 5466 16836 5488
rect 1104 5414 4898 5466
rect 4950 5414 4962 5466
rect 5014 5414 5026 5466
rect 5078 5414 5090 5466
rect 5142 5414 5154 5466
rect 5206 5414 8846 5466
rect 8898 5414 8910 5466
rect 8962 5414 8974 5466
rect 9026 5414 9038 5466
rect 9090 5414 9102 5466
rect 9154 5414 12794 5466
rect 12846 5414 12858 5466
rect 12910 5414 12922 5466
rect 12974 5414 12986 5466
rect 13038 5414 13050 5466
rect 13102 5414 16836 5466
rect 1104 5392 16836 5414
rect 1946 5312 1952 5364
rect 2004 5352 2010 5364
rect 2590 5352 2596 5364
rect 2004 5324 2596 5352
rect 2004 5312 2010 5324
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 6454 5352 6460 5364
rect 3988 5324 6460 5352
rect 842 5244 848 5296
rect 900 5284 906 5296
rect 3988 5284 4016 5324
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6546 5312 6552 5364
rect 6604 5312 6610 5364
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 9217 5355 9275 5361
rect 9217 5352 9229 5355
rect 7892 5324 9229 5352
rect 7892 5312 7898 5324
rect 9217 5321 9229 5324
rect 9263 5321 9275 5355
rect 10778 5352 10784 5364
rect 9217 5315 9275 5321
rect 9784 5324 10784 5352
rect 6270 5284 6276 5296
rect 900 5256 1992 5284
rect 900 5244 906 5256
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5176 1458 5228
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 1854 5216 1860 5228
rect 1719 5188 1860 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 1762 5148 1768 5160
rect 1723 5120 1768 5148
rect 1762 5108 1768 5120
rect 1820 5108 1826 5160
rect 1964 5148 1992 5256
rect 2240 5256 4016 5284
rect 5184 5256 6276 5284
rect 2240 5225 2268 5256
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5185 2283 5219
rect 2481 5219 2539 5225
rect 2481 5216 2493 5219
rect 2225 5179 2283 5185
rect 2332 5188 2493 5216
rect 2332 5148 2360 5188
rect 2481 5185 2493 5188
rect 2527 5185 2539 5219
rect 2481 5179 2539 5185
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5216 4123 5219
rect 5074 5216 5080 5228
rect 4111 5188 5080 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 1964 5120 2360 5148
rect 3326 5108 3332 5160
rect 3384 5148 3390 5160
rect 3694 5148 3700 5160
rect 3384 5120 3700 5148
rect 3384 5108 3390 5120
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 5184 5080 5212 5256
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 6564 5231 6592 5312
rect 7006 5284 7012 5296
rect 6886 5256 7012 5284
rect 6553 5225 6611 5231
rect 6886 5225 6914 5256
rect 7006 5244 7012 5256
rect 7064 5244 7070 5296
rect 7926 5244 7932 5296
rect 7984 5284 7990 5296
rect 7984 5256 8029 5284
rect 7984 5244 7990 5256
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 3160 5052 5212 5080
rect 6104 5188 6377 5216
rect 2590 4972 2596 5024
rect 2648 5012 2654 5024
rect 3160 5012 3188 5052
rect 2648 4984 3188 5012
rect 3605 5015 3663 5021
rect 2648 4972 2654 4984
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 5166 5012 5172 5024
rect 3651 4984 5172 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 5350 5012 5356 5024
rect 5311 4984 5356 5012
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 6104 5012 6132 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6553 5191 6565 5225
rect 6599 5191 6611 5225
rect 6553 5185 6611 5191
rect 6872 5219 6930 5225
rect 6872 5185 6884 5219
rect 6918 5185 6930 5219
rect 9122 5216 9128 5228
rect 6365 5179 6423 5185
rect 6872 5179 6930 5185
rect 7024 5188 9128 5216
rect 6638 5148 6644 5160
rect 6599 5120 6644 5148
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5148 6791 5151
rect 7024 5148 7052 5188
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 6779 5120 7052 5148
rect 7101 5151 7159 5157
rect 6779 5117 6791 5120
rect 6733 5111 6791 5117
rect 7101 5117 7113 5151
rect 7147 5148 7159 5151
rect 9784 5148 9812 5324
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 11517 5355 11575 5361
rect 11517 5321 11529 5355
rect 11563 5352 11575 5355
rect 15470 5352 15476 5364
rect 11563 5324 15476 5352
rect 11563 5321 11575 5324
rect 11517 5315 11575 5321
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 9858 5244 9864 5296
rect 9916 5284 9922 5296
rect 9916 5256 10088 5284
rect 9916 5244 9922 5256
rect 7147 5120 9812 5148
rect 10060 5148 10088 5256
rect 10686 5244 10692 5296
rect 10744 5284 10750 5296
rect 11885 5287 11943 5293
rect 10744 5256 11744 5284
rect 10744 5244 10750 5256
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 10060 5120 10149 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 10226 5108 10232 5160
rect 10284 5148 10290 5160
rect 10336 5148 10364 5179
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 10560 5188 10609 5216
rect 10560 5176 10566 5188
rect 10597 5185 10609 5188
rect 10643 5216 10655 5219
rect 11238 5216 11244 5228
rect 10643 5188 11244 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 11238 5176 11244 5188
rect 11296 5176 11302 5228
rect 11716 5225 11744 5256
rect 11885 5253 11897 5287
rect 11931 5284 11943 5287
rect 12526 5284 12532 5296
rect 11931 5256 12532 5284
rect 11931 5253 11943 5256
rect 11885 5247 11943 5253
rect 12526 5244 12532 5256
rect 12584 5244 12590 5296
rect 12805 5287 12863 5293
rect 12805 5253 12817 5287
rect 12851 5284 12863 5287
rect 13170 5284 13176 5296
rect 12851 5256 13176 5284
rect 12851 5253 12863 5256
rect 12805 5247 12863 5253
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 13446 5244 13452 5296
rect 13504 5284 13510 5296
rect 15349 5287 15407 5293
rect 15349 5284 15361 5287
rect 13504 5256 15361 5284
rect 13504 5244 13510 5256
rect 15349 5253 15361 5256
rect 15395 5253 15407 5287
rect 15349 5247 15407 5253
rect 15565 5287 15623 5293
rect 15565 5253 15577 5287
rect 15611 5284 15623 5287
rect 15611 5256 15976 5284
rect 15611 5253 15623 5256
rect 15565 5247 15623 5253
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11974 5216 11980 5228
rect 11935 5188 11980 5216
rect 11701 5179 11759 5185
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 12158 5176 12164 5228
rect 12216 5216 12222 5228
rect 12342 5216 12348 5228
rect 12216 5188 12348 5216
rect 12216 5176 12222 5188
rect 12342 5176 12348 5188
rect 12400 5176 12406 5228
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 13354 5216 13360 5228
rect 12492 5188 13360 5216
rect 12492 5176 12498 5188
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 14553 5219 14611 5225
rect 14553 5185 14565 5219
rect 14599 5216 14611 5219
rect 15838 5216 15844 5228
rect 14599 5188 15844 5216
rect 14599 5185 14611 5188
rect 14553 5179 14611 5185
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 10284 5120 10364 5148
rect 10413 5151 10471 5157
rect 10284 5108 10290 5120
rect 10413 5117 10425 5151
rect 10459 5148 10471 5151
rect 10459 5120 10732 5148
rect 10459 5117 10471 5120
rect 10413 5111 10471 5117
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 9858 5080 9864 5092
rect 6880 5052 9864 5080
rect 6880 5040 6886 5052
rect 9858 5040 9864 5052
rect 9916 5040 9922 5092
rect 9950 5040 9956 5092
rect 10008 5080 10014 5092
rect 10318 5080 10324 5092
rect 10008 5052 10324 5080
rect 10008 5040 10014 5052
rect 10318 5040 10324 5052
rect 10376 5040 10382 5092
rect 10505 5083 10563 5089
rect 10505 5049 10517 5083
rect 10551 5080 10563 5083
rect 10594 5080 10600 5092
rect 10551 5052 10600 5080
rect 10551 5049 10563 5052
rect 10505 5043 10563 5049
rect 10594 5040 10600 5052
rect 10652 5040 10658 5092
rect 10704 5080 10732 5120
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 13998 5148 14004 5160
rect 10836 5120 14004 5148
rect 10836 5108 10842 5120
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 15948 5148 15976 5256
rect 14844 5120 15976 5148
rect 11882 5080 11888 5092
rect 10704 5052 11888 5080
rect 11882 5040 11888 5052
rect 11940 5040 11946 5092
rect 12342 5080 12348 5092
rect 12176 5052 12348 5080
rect 8662 5012 8668 5024
rect 6104 4984 8668 5012
rect 8662 4972 8668 4984
rect 8720 4972 8726 5024
rect 8938 4972 8944 5024
rect 8996 5012 9002 5024
rect 12176 5012 12204 5052
rect 12342 5040 12348 5052
rect 12400 5040 12406 5092
rect 12802 5040 12808 5092
rect 12860 5080 12866 5092
rect 14844 5089 14872 5120
rect 14829 5083 14887 5089
rect 14829 5080 14841 5083
rect 12860 5052 14841 5080
rect 12860 5040 12866 5052
rect 14829 5049 14841 5052
rect 14875 5049 14887 5083
rect 14829 5043 14887 5049
rect 8996 4984 12204 5012
rect 8996 4972 9002 4984
rect 12250 4972 12256 5024
rect 12308 5012 12314 5024
rect 12894 5012 12900 5024
rect 12308 4984 12900 5012
rect 12308 4972 12314 4984
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 12986 4972 12992 5024
rect 13044 5012 13050 5024
rect 14274 5012 14280 5024
rect 13044 4984 14280 5012
rect 13044 4972 13050 4984
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 15194 5012 15200 5024
rect 15155 4984 15200 5012
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15286 4972 15292 5024
rect 15344 5012 15350 5024
rect 15381 5015 15439 5021
rect 15381 5012 15393 5015
rect 15344 4984 15393 5012
rect 15344 4972 15350 4984
rect 15381 4981 15393 4984
rect 15427 5012 15439 5015
rect 15470 5012 15476 5024
rect 15427 4984 15476 5012
rect 15427 4981 15439 4984
rect 15381 4975 15439 4981
rect 15470 4972 15476 4984
rect 15528 4972 15534 5024
rect 1104 4922 16836 4944
rect 1104 4870 2924 4922
rect 2976 4870 2988 4922
rect 3040 4870 3052 4922
rect 3104 4870 3116 4922
rect 3168 4870 3180 4922
rect 3232 4870 6872 4922
rect 6924 4870 6936 4922
rect 6988 4870 7000 4922
rect 7052 4870 7064 4922
rect 7116 4870 7128 4922
rect 7180 4870 10820 4922
rect 10872 4870 10884 4922
rect 10936 4870 10948 4922
rect 11000 4870 11012 4922
rect 11064 4870 11076 4922
rect 11128 4870 14768 4922
rect 14820 4870 14832 4922
rect 14884 4870 14896 4922
rect 14948 4870 14960 4922
rect 15012 4870 15024 4922
rect 15076 4870 16836 4922
rect 1104 4848 16836 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 3142 4808 3148 4820
rect 1820 4780 3148 4808
rect 1820 4768 1826 4780
rect 3142 4768 3148 4780
rect 3200 4808 3206 4820
rect 3786 4808 3792 4820
rect 3200 4780 3792 4808
rect 3200 4768 3206 4780
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4246 4808 4252 4820
rect 3988 4780 4252 4808
rect 2590 4740 2596 4752
rect 2551 4712 2596 4740
rect 2590 4700 2596 4712
rect 2648 4700 2654 4752
rect 3988 4740 4016 4780
rect 4246 4768 4252 4780
rect 4304 4768 4310 4820
rect 5074 4768 5080 4820
rect 5132 4808 5138 4820
rect 7834 4808 7840 4820
rect 5132 4780 7840 4808
rect 5132 4768 5138 4780
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 8220 4780 9812 4808
rect 2700 4712 4016 4740
rect 1486 4672 1492 4684
rect 1447 4644 1492 4672
rect 1486 4632 1492 4644
rect 1544 4632 1550 4684
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 1596 4536 1624 4567
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 2222 4604 2228 4616
rect 1820 4576 2228 4604
rect 1820 4564 1826 4576
rect 2222 4564 2228 4576
rect 2280 4564 2286 4616
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 2700 4613 2728 4712
rect 4062 4700 4068 4752
rect 4120 4700 4126 4752
rect 8220 4740 8248 4780
rect 7668 4712 8248 4740
rect 3234 4672 3240 4684
rect 2884 4644 3240 4672
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 2884 4536 2912 4644
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 4080 4672 4108 4700
rect 7668 4672 7696 4712
rect 8294 4700 8300 4752
rect 8352 4740 8358 4752
rect 8938 4740 8944 4752
rect 8352 4712 8397 4740
rect 8899 4712 8944 4740
rect 8352 4700 8358 4712
rect 8938 4700 8944 4712
rect 8996 4700 9002 4752
rect 9122 4700 9128 4752
rect 9180 4740 9186 4752
rect 9784 4740 9812 4780
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 12066 4808 12072 4820
rect 9916 4780 12072 4808
rect 9916 4768 9922 4780
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12621 4811 12679 4817
rect 12621 4808 12633 4811
rect 12360 4780 12633 4808
rect 12360 4752 12388 4780
rect 12621 4777 12633 4780
rect 12667 4777 12679 4811
rect 12986 4808 12992 4820
rect 12947 4780 12992 4808
rect 12621 4771 12679 4777
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 14274 4808 14280 4820
rect 14235 4780 14280 4808
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 15841 4811 15899 4817
rect 15841 4808 15853 4811
rect 14384 4780 15853 4808
rect 10410 4740 10416 4752
rect 9180 4712 9625 4740
rect 9784 4712 10416 4740
rect 9180 4700 9186 4712
rect 3436 4644 4108 4672
rect 5276 4644 7696 4672
rect 7929 4675 7987 4681
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4573 3019 4607
rect 3142 4604 3148 4616
rect 3103 4576 3148 4604
rect 2961 4567 3019 4573
rect 1596 4508 2912 4536
rect 2976 4536 3004 4567
rect 3142 4564 3148 4576
rect 3200 4604 3206 4616
rect 3326 4604 3332 4616
rect 3200 4576 3332 4604
rect 3200 4564 3206 4576
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 3436 4536 3464 4644
rect 3786 4604 3792 4616
rect 3747 4576 3792 4604
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 4062 4604 4068 4616
rect 4023 4576 4068 4604
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 5276 4613 5304 4644
rect 7929 4641 7941 4675
rect 7975 4672 7987 4675
rect 8018 4672 8024 4684
rect 7975 4644 8024 4672
rect 7975 4641 7987 4644
rect 7929 4635 7987 4641
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 8662 4672 8668 4684
rect 8220 4644 8668 4672
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 8220 4604 8248 4644
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 9401 4675 9459 4681
rect 9401 4641 9413 4675
rect 9447 4672 9459 4675
rect 9490 4672 9496 4684
rect 9447 4644 9496 4672
rect 9447 4641 9459 4644
rect 9401 4635 9459 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 9597 4672 9625 4712
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 12342 4700 12348 4752
rect 12400 4700 12406 4752
rect 12802 4700 12808 4752
rect 12860 4740 12866 4752
rect 14384 4740 14412 4780
rect 15841 4777 15853 4780
rect 15887 4777 15899 4811
rect 15841 4771 15899 4777
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 15988 4780 16033 4808
rect 15988 4768 15994 4780
rect 12860 4712 14412 4740
rect 12860 4700 12866 4712
rect 14918 4700 14924 4752
rect 14976 4740 14982 4752
rect 15013 4743 15071 4749
rect 15013 4740 15025 4743
rect 14976 4712 15025 4740
rect 14976 4700 14982 4712
rect 15013 4709 15025 4712
rect 15059 4709 15071 4743
rect 15013 4703 15071 4709
rect 12526 4672 12532 4684
rect 9597 4644 12532 4672
rect 12526 4632 12532 4644
rect 12584 4672 12590 4684
rect 12713 4675 12771 4681
rect 12713 4672 12725 4675
rect 12584 4644 12725 4672
rect 12584 4632 12590 4644
rect 12713 4641 12725 4644
rect 12759 4672 12771 4675
rect 16025 4675 16083 4681
rect 16025 4672 16037 4675
rect 12759 4644 16037 4672
rect 12759 4641 12771 4644
rect 12713 4635 12771 4641
rect 16025 4641 16037 4644
rect 16071 4641 16083 4675
rect 16025 4635 16083 4641
rect 9122 4604 9128 4616
rect 7055 4576 7788 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 2976 4508 3464 4536
rect 5810 4496 5816 4548
rect 5868 4536 5874 4548
rect 6546 4536 6552 4548
rect 5868 4508 6552 4536
rect 5868 4496 5874 4508
rect 6546 4496 6552 4508
rect 6604 4496 6610 4548
rect 7760 4536 7788 4576
rect 8036 4576 8248 4604
rect 9083 4576 9128 4604
rect 8036 4536 8064 4576
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4604 9367 4607
rect 10226 4604 10232 4616
rect 9355 4576 10232 4604
rect 9355 4573 9367 4576
rect 9309 4567 9367 4573
rect 9232 4536 9260 4567
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4604 10471 4607
rect 10778 4604 10784 4616
rect 10459 4576 10784 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 10778 4564 10784 4576
rect 10836 4564 10842 4616
rect 10962 4564 10968 4616
rect 11020 4604 11026 4616
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 11020 4576 12633 4604
rect 11020 4564 11026 4576
rect 12621 4573 12633 4576
rect 12667 4604 12679 4607
rect 12802 4604 12808 4616
rect 12667 4576 12808 4604
rect 12667 4573 12679 4576
rect 12621 4567 12679 4573
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 14921 4607 14979 4613
rect 14921 4604 14933 4607
rect 13412 4576 14933 4604
rect 13412 4564 13418 4576
rect 14921 4573 14933 4576
rect 14967 4573 14979 4607
rect 14921 4567 14979 4573
rect 15105 4607 15163 4613
rect 15105 4573 15117 4607
rect 15151 4573 15163 4607
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15105 4567 15163 4573
rect 15212 4576 15761 4604
rect 7760 4508 8064 4536
rect 8128 4508 9260 4536
rect 1949 4471 2007 4477
rect 1949 4437 1961 4471
rect 1995 4468 2007 4471
rect 6730 4468 6736 4480
rect 1995 4440 6736 4468
rect 1995 4437 2007 4440
rect 1949 4431 2007 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 8018 4428 8024 4480
rect 8076 4468 8082 4480
rect 8128 4468 8156 4508
rect 9766 4496 9772 4548
rect 9824 4536 9830 4548
rect 12161 4539 12219 4545
rect 9824 4508 11376 4536
rect 9824 4496 9830 4508
rect 8076 4440 8156 4468
rect 8389 4471 8447 4477
rect 8076 4428 8082 4440
rect 8389 4437 8401 4471
rect 8435 4468 8447 4471
rect 8846 4468 8852 4480
rect 8435 4440 8852 4468
rect 8435 4437 8447 4440
rect 8389 4431 8447 4437
rect 8846 4428 8852 4440
rect 8904 4428 8910 4480
rect 9122 4428 9128 4480
rect 9180 4468 9186 4480
rect 11238 4468 11244 4480
rect 9180 4440 11244 4468
rect 9180 4428 9186 4440
rect 11238 4428 11244 4440
rect 11296 4428 11302 4480
rect 11348 4468 11376 4508
rect 12161 4505 12173 4539
rect 12207 4536 12219 4539
rect 12250 4536 12256 4548
rect 12207 4508 12256 4536
rect 12207 4505 12219 4508
rect 12161 4499 12219 4505
rect 12250 4496 12256 4508
rect 12308 4496 12314 4548
rect 12894 4496 12900 4548
rect 12952 4536 12958 4548
rect 14093 4539 14151 4545
rect 14093 4536 14105 4539
rect 12952 4508 14105 4536
rect 12952 4496 12958 4508
rect 14093 4505 14105 4508
rect 14139 4505 14151 4539
rect 14093 4499 14151 4505
rect 14309 4539 14367 4545
rect 14309 4505 14321 4539
rect 14355 4536 14367 4539
rect 14642 4536 14648 4548
rect 14355 4508 14648 4536
rect 14355 4505 14367 4508
rect 14309 4499 14367 4505
rect 14642 4496 14648 4508
rect 14700 4496 14706 4548
rect 14734 4496 14740 4548
rect 14792 4536 14798 4548
rect 15120 4536 15148 4567
rect 14792 4508 15148 4536
rect 14792 4496 14798 4508
rect 13446 4468 13452 4480
rect 11348 4440 13452 4468
rect 13446 4428 13452 4440
rect 13504 4428 13510 4480
rect 14458 4468 14464 4480
rect 14419 4440 14464 4468
rect 14458 4428 14464 4440
rect 14516 4468 14522 4480
rect 15212 4468 15240 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 14516 4440 15240 4468
rect 14516 4428 14522 4440
rect 1104 4378 16836 4400
rect 1104 4326 4898 4378
rect 4950 4326 4962 4378
rect 5014 4326 5026 4378
rect 5078 4326 5090 4378
rect 5142 4326 5154 4378
rect 5206 4326 8846 4378
rect 8898 4326 8910 4378
rect 8962 4326 8974 4378
rect 9026 4326 9038 4378
rect 9090 4326 9102 4378
rect 9154 4326 12794 4378
rect 12846 4326 12858 4378
rect 12910 4326 12922 4378
rect 12974 4326 12986 4378
rect 13038 4326 13050 4378
rect 13102 4326 16836 4378
rect 1104 4304 16836 4326
rect 2498 4264 2504 4276
rect 1412 4236 2504 4264
rect 1412 4137 1440 4236
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 6454 4224 6460 4276
rect 6512 4264 6518 4276
rect 9490 4264 9496 4276
rect 6512 4236 9496 4264
rect 6512 4224 6518 4236
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 10962 4264 10968 4276
rect 9824 4236 10968 4264
rect 9824 4224 9830 4236
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 11054 4224 11060 4276
rect 11112 4264 11118 4276
rect 11885 4267 11943 4273
rect 11885 4264 11897 4267
rect 11112 4236 11897 4264
rect 11112 4224 11118 4236
rect 11885 4233 11897 4236
rect 11931 4233 11943 4267
rect 11885 4227 11943 4233
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 14458 4264 14464 4276
rect 12492 4236 14464 4264
rect 12492 4224 12498 4236
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 14826 4224 14832 4276
rect 14884 4264 14890 4276
rect 16758 4264 16764 4276
rect 14884 4236 16764 4264
rect 14884 4224 14890 4236
rect 16758 4224 16764 4236
rect 16816 4224 16822 4276
rect 1765 4199 1823 4205
rect 1765 4165 1777 4199
rect 1811 4196 1823 4199
rect 1946 4196 1952 4208
rect 1811 4168 1952 4196
rect 1811 4165 1823 4168
rect 1765 4159 1823 4165
rect 1946 4156 1952 4168
rect 2004 4196 2010 4208
rect 2406 4196 2412 4208
rect 2004 4168 2412 4196
rect 2004 4156 2010 4168
rect 2406 4156 2412 4168
rect 2464 4156 2470 4208
rect 2866 4205 2872 4208
rect 2860 4196 2872 4205
rect 2827 4168 2872 4196
rect 2860 4159 2872 4168
rect 2866 4156 2872 4159
rect 2924 4156 2930 4208
rect 2976 4168 6592 4196
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 2498 4088 2504 4140
rect 2556 4128 2562 4140
rect 2976 4128 3004 4168
rect 4430 4128 4436 4140
rect 2556 4100 3004 4128
rect 4391 4100 4436 4128
rect 2556 4088 2562 4100
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 6564 4137 6592 4168
rect 7024 4168 7512 4196
rect 4689 4131 4747 4137
rect 4689 4128 4701 4131
rect 4540 4100 4701 4128
rect 658 4020 664 4072
rect 716 4060 722 4072
rect 2590 4060 2596 4072
rect 716 4032 2452 4060
rect 2551 4032 2596 4060
rect 716 4020 722 4032
rect 2222 3992 2228 4004
rect 1780 3964 2228 3992
rect 1780 3933 1808 3964
rect 2222 3952 2228 3964
rect 2280 3952 2286 4004
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3893 1823 3927
rect 1765 3887 1823 3893
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3924 2007 3927
rect 2314 3924 2320 3936
rect 1995 3896 2320 3924
rect 1995 3893 2007 3896
rect 1949 3887 2007 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2424 3924 2452 4032
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 4540 4060 4568 4100
rect 4689 4097 4701 4100
rect 4735 4097 4747 4131
rect 4689 4091 4747 4097
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 6914 4128 6920 4140
rect 6595 4100 6920 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 6822 4060 6828 4072
rect 3712 4032 4568 4060
rect 5828 4032 6828 4060
rect 3712 3924 3740 4032
rect 3786 3952 3792 4004
rect 3844 3992 3850 4004
rect 3973 3995 4031 4001
rect 3973 3992 3985 3995
rect 3844 3964 3985 3992
rect 3844 3952 3850 3964
rect 3973 3961 3985 3964
rect 4019 3961 4031 3995
rect 3973 3955 4031 3961
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 5718 3992 5724 4004
rect 5592 3964 5724 3992
rect 5592 3952 5598 3964
rect 5718 3952 5724 3964
rect 5776 3952 5782 4004
rect 5828 4001 5856 4032
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 5813 3995 5871 4001
rect 5813 3961 5825 3995
rect 5859 3961 5871 3995
rect 6362 3992 6368 4004
rect 6323 3964 6368 3992
rect 5813 3955 5871 3961
rect 6362 3952 6368 3964
rect 6420 3952 6426 4004
rect 7024 3992 7052 4168
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7190 4128 7196 4140
rect 7147 4100 7196 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 7374 4137 7380 4140
rect 7368 4128 7380 4137
rect 7335 4100 7380 4128
rect 7368 4091 7380 4100
rect 7374 4088 7380 4091
rect 7432 4088 7438 4140
rect 7484 4128 7512 4168
rect 8662 4156 8668 4208
rect 8720 4196 8726 4208
rect 8938 4196 8944 4208
rect 8720 4168 8944 4196
rect 8720 4156 8726 4168
rect 8938 4156 8944 4168
rect 8996 4196 9002 4208
rect 11514 4196 11520 4208
rect 8996 4168 11520 4196
rect 8996 4156 9002 4168
rect 11514 4156 11520 4168
rect 11572 4156 11578 4208
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 11664 4168 11744 4196
rect 11664 4156 11670 4168
rect 8846 4128 8852 4140
rect 7484 4100 8852 4128
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 9214 4128 9220 4140
rect 9175 4100 9220 4128
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 9674 4088 9680 4140
rect 9732 4128 9738 4140
rect 11716 4137 11744 4168
rect 11790 4156 11796 4208
rect 11848 4196 11854 4208
rect 12158 4196 12164 4208
rect 11848 4168 12164 4196
rect 11848 4156 11854 4168
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 12250 4156 12256 4208
rect 12308 4196 12314 4208
rect 13262 4196 13268 4208
rect 12308 4168 13268 4196
rect 12308 4156 12314 4168
rect 11701 4131 11759 4137
rect 9732 4100 11652 4128
rect 9732 4088 9738 4100
rect 8478 4020 8484 4072
rect 8536 4060 8542 4072
rect 8662 4060 8668 4072
rect 8536 4032 8668 4060
rect 8536 4020 8542 4032
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 9766 4060 9772 4072
rect 9548 4032 9772 4060
rect 9548 4020 9554 4032
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 10778 4060 10784 4072
rect 10652 4032 10784 4060
rect 10652 4020 10658 4032
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 11204 4032 11529 4060
rect 11204 4020 11210 4032
rect 11517 4029 11529 4032
rect 11563 4029 11575 4063
rect 11624 4060 11652 4100
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 11992 4060 12020 4091
rect 12066 4088 12072 4140
rect 12124 4128 12130 4140
rect 12342 4128 12348 4140
rect 12124 4100 12348 4128
rect 12124 4088 12130 4100
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 13096 4137 13124 4168
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 13722 4156 13728 4208
rect 13780 4196 13786 4208
rect 14918 4196 14924 4208
rect 13780 4168 14924 4196
rect 13780 4156 13786 4168
rect 14918 4156 14924 4168
rect 14976 4156 14982 4208
rect 15930 4156 15936 4208
rect 15988 4196 15994 4208
rect 15988 4168 16160 4196
rect 15988 4156 15994 4168
rect 13081 4131 13139 4137
rect 13081 4097 13093 4131
rect 13127 4097 13139 4131
rect 13081 4091 13139 4097
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13219 4100 13492 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 13464 4072 13492 4100
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13596 4100 13829 4128
rect 13596 4088 13602 4100
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 14090 4128 14096 4140
rect 14051 4100 14096 4128
rect 13817 4091 13875 4097
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 14737 4131 14795 4137
rect 14737 4128 14749 4131
rect 14516 4100 14749 4128
rect 14516 4088 14522 4100
rect 14737 4097 14749 4100
rect 14783 4128 14795 4131
rect 14826 4128 14832 4140
rect 14783 4100 14832 4128
rect 14783 4097 14795 4100
rect 14737 4091 14795 4097
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 16022 4128 16028 4140
rect 15983 4100 16028 4128
rect 15841 4091 15899 4097
rect 11624 4032 12020 4060
rect 11517 4023 11575 4029
rect 12158 4020 12164 4072
rect 12216 4060 12222 4072
rect 13357 4063 13415 4069
rect 13357 4060 13369 4063
rect 12216 4032 13369 4060
rect 12216 4020 12222 4032
rect 13357 4029 13369 4032
rect 13403 4029 13415 4063
rect 13357 4023 13415 4029
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 13504 4032 14044 4060
rect 13504 4020 13510 4032
rect 6472 3964 7052 3992
rect 2424 3896 3740 3924
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6472 3924 6500 3964
rect 8202 3952 8208 4004
rect 8260 3992 8266 4004
rect 13909 3995 13967 4001
rect 13909 3992 13921 3995
rect 8260 3964 12434 3992
rect 8260 3952 8266 3964
rect 6144 3896 6500 3924
rect 6144 3884 6150 3896
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 8294 3924 8300 3936
rect 6696 3896 8300 3924
rect 6696 3884 6702 3896
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8478 3924 8484 3936
rect 8439 3896 8484 3924
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 8846 3884 8852 3936
rect 8904 3924 8910 3936
rect 12250 3924 12256 3936
rect 8904 3896 12256 3924
rect 8904 3884 8910 3896
rect 12250 3884 12256 3896
rect 12308 3884 12314 3936
rect 12406 3924 12434 3964
rect 13004 3964 13921 3992
rect 13004 3924 13032 3964
rect 13909 3961 13921 3964
rect 13955 3961 13967 3995
rect 14016 3992 14044 4032
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14921 4063 14979 4069
rect 14921 4060 14933 4063
rect 14424 4032 14933 4060
rect 14424 4020 14430 4032
rect 14921 4029 14933 4032
rect 14967 4029 14979 4063
rect 14921 4023 14979 4029
rect 15102 4020 15108 4072
rect 15160 4060 15166 4072
rect 15856 4060 15884 4091
rect 16022 4088 16028 4100
rect 16080 4088 16086 4140
rect 16132 4137 16160 4168
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 16850 4060 16856 4072
rect 15160 4032 16856 4060
rect 15160 4020 15166 4032
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 14734 3992 14740 4004
rect 14016 3964 14740 3992
rect 13909 3955 13967 3961
rect 14734 3952 14740 3964
rect 14792 3952 14798 4004
rect 12406 3896 13032 3924
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 14550 3924 14556 3936
rect 14332 3896 14556 3924
rect 14332 3884 14338 3896
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 15286 3884 15292 3936
rect 15344 3924 15350 3936
rect 15841 3927 15899 3933
rect 15841 3924 15853 3927
rect 15344 3896 15853 3924
rect 15344 3884 15350 3896
rect 15841 3893 15853 3896
rect 15887 3893 15899 3927
rect 15841 3887 15899 3893
rect 1104 3834 16836 3856
rect 1104 3782 2924 3834
rect 2976 3782 2988 3834
rect 3040 3782 3052 3834
rect 3104 3782 3116 3834
rect 3168 3782 3180 3834
rect 3232 3782 6872 3834
rect 6924 3782 6936 3834
rect 6988 3782 7000 3834
rect 7052 3782 7064 3834
rect 7116 3782 7128 3834
rect 7180 3782 10820 3834
rect 10872 3782 10884 3834
rect 10936 3782 10948 3834
rect 11000 3782 11012 3834
rect 11064 3782 11076 3834
rect 11128 3782 14768 3834
rect 14820 3782 14832 3834
rect 14884 3782 14896 3834
rect 14948 3782 14960 3834
rect 15012 3782 15024 3834
rect 15076 3782 16836 3834
rect 1104 3760 16836 3782
rect 3510 3720 3516 3732
rect 1780 3692 3516 3720
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 1780 3584 1808 3692
rect 3510 3680 3516 3692
rect 3568 3720 3574 3732
rect 6086 3720 6092 3732
rect 3568 3692 6092 3720
rect 3568 3680 3574 3692
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 6638 3720 6644 3732
rect 6236 3692 6644 3720
rect 6236 3680 6242 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 6733 3723 6791 3729
rect 6733 3689 6745 3723
rect 6779 3720 6791 3723
rect 7098 3720 7104 3732
rect 6779 3692 7104 3720
rect 6779 3689 6791 3692
rect 6733 3683 6791 3689
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 10962 3720 10968 3732
rect 7300 3692 9996 3720
rect 10923 3692 10968 3720
rect 2961 3655 3019 3661
rect 2961 3621 2973 3655
rect 3007 3621 3019 3655
rect 2961 3615 3019 3621
rect 1719 3556 1808 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 1946 3544 1952 3596
rect 2004 3584 2010 3596
rect 2498 3584 2504 3596
rect 2004 3556 2504 3584
rect 2004 3544 2010 3556
rect 2498 3544 2504 3556
rect 2556 3544 2562 3596
rect 2976 3584 3004 3615
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 4706 3652 4712 3664
rect 4212 3624 4712 3652
rect 4212 3612 4218 3624
rect 4706 3612 4712 3624
rect 4764 3612 4770 3664
rect 7190 3652 7196 3664
rect 5184 3624 7196 3652
rect 4065 3587 4123 3593
rect 2976 3556 4016 3584
rect 3142 3516 3148 3528
rect 3103 3488 3148 3516
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3326 3516 3332 3528
rect 3283 3488 3332 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3326 3476 3332 3488
rect 3384 3516 3390 3528
rect 3510 3516 3516 3528
rect 3384 3488 3516 3516
rect 3384 3476 3390 3488
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 3786 3516 3792 3528
rect 3747 3488 3792 3516
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 3988 3516 4016 3556
rect 4065 3553 4077 3587
rect 4111 3584 4123 3587
rect 4246 3584 4252 3596
rect 4111 3556 4252 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 4246 3544 4252 3556
rect 4304 3584 4310 3596
rect 4522 3584 4528 3596
rect 4304 3556 4528 3584
rect 4304 3544 4310 3556
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 5184 3516 5212 3624
rect 7190 3612 7196 3624
rect 7248 3612 7254 3664
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 7300 3584 7328 3692
rect 9968 3664 9996 3692
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 12250 3720 12256 3732
rect 11940 3692 12256 3720
rect 11940 3680 11946 3692
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 12342 3680 12348 3732
rect 12400 3720 12406 3732
rect 13173 3723 13231 3729
rect 13173 3720 13185 3723
rect 12400 3692 13185 3720
rect 12400 3680 12406 3692
rect 13173 3689 13185 3692
rect 13219 3689 13231 3723
rect 14274 3720 14280 3732
rect 14235 3692 14280 3720
rect 13173 3683 13231 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 16482 3720 16488 3732
rect 14608 3692 16488 3720
rect 14608 3680 14614 3692
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 8018 3652 8024 3664
rect 7979 3624 8024 3652
rect 8018 3612 8024 3624
rect 8076 3612 8082 3664
rect 9950 3612 9956 3664
rect 10008 3612 10014 3664
rect 11698 3652 11704 3664
rect 11659 3624 11704 3652
rect 11698 3612 11704 3624
rect 11756 3612 11762 3664
rect 12158 3612 12164 3664
rect 12216 3652 12222 3664
rect 14292 3652 14320 3680
rect 12216 3624 14320 3652
rect 15473 3655 15531 3661
rect 12216 3612 12222 3624
rect 15473 3621 15485 3655
rect 15519 3652 15531 3655
rect 15746 3652 15752 3664
rect 15519 3624 15752 3652
rect 15519 3621 15531 3624
rect 15473 3615 15531 3621
rect 15746 3612 15752 3624
rect 15804 3612 15810 3664
rect 8938 3584 8944 3596
rect 6604 3556 7604 3584
rect 8899 3556 8944 3584
rect 6604 3544 6610 3556
rect 3988 3488 5212 3516
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 5442 3516 5448 3528
rect 5307 3488 5448 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 7282 3516 7288 3528
rect 6512 3488 7288 3516
rect 6512 3476 6518 3488
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 7576 3510 7604 3556
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 10284 3556 10824 3584
rect 10284 3544 10290 3556
rect 7653 3519 7711 3525
rect 7653 3510 7665 3519
rect 7576 3485 7665 3510
rect 7699 3485 7711 3519
rect 7576 3482 7711 3485
rect 7653 3479 7711 3482
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3516 7895 3519
rect 7883 3488 7972 3516
rect 7883 3485 7895 3488
rect 7837 3479 7895 3485
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 2961 3451 3019 3457
rect 2961 3448 2973 3451
rect 992 3420 2973 3448
rect 992 3408 998 3420
rect 2961 3417 2973 3420
rect 3007 3417 3019 3451
rect 2961 3411 3019 3417
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 6178 3448 6184 3460
rect 3752 3420 6184 3448
rect 3752 3408 3758 3420
rect 6178 3408 6184 3420
rect 6236 3408 6242 3460
rect 7374 3448 7380 3460
rect 6288 3420 7380 3448
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 6288 3380 6316 3420
rect 7374 3408 7380 3420
rect 7432 3408 7438 3460
rect 7484 3448 7512 3479
rect 7742 3448 7748 3460
rect 7484 3420 7604 3448
rect 7655 3420 7748 3448
rect 7576 3392 7604 3420
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 7944 3448 7972 3488
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 9197 3519 9255 3525
rect 9197 3516 9209 3519
rect 8168 3488 9209 3516
rect 8168 3476 8174 3488
rect 9197 3485 9209 3488
rect 9243 3485 9255 3519
rect 9197 3479 9255 3485
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 9968 3516 10180 3518
rect 10796 3516 10824 3556
rect 11054 3544 11060 3596
rect 11112 3584 11118 3596
rect 14921 3587 14979 3593
rect 14921 3584 14933 3587
rect 11112 3556 14933 3584
rect 11112 3544 11118 3556
rect 14921 3553 14933 3556
rect 14967 3553 14979 3587
rect 14921 3547 14979 3553
rect 11238 3516 11244 3528
rect 9548 3492 10548 3516
rect 9548 3490 10640 3492
rect 9548 3488 9996 3490
rect 10152 3488 10640 3490
rect 9548 3476 9554 3488
rect 10520 3464 10640 3488
rect 8202 3448 8208 3460
rect 7944 3420 8208 3448
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 2924 3352 6316 3380
rect 2924 3340 2930 3352
rect 7558 3340 7564 3392
rect 7616 3340 7622 3392
rect 7760 3380 7788 3408
rect 10321 3383 10379 3389
rect 10321 3380 10333 3383
rect 7760 3352 10333 3380
rect 10321 3349 10333 3352
rect 10367 3349 10379 3383
rect 10612 3380 10640 3464
rect 10796 3488 11244 3516
rect 10796 3460 10824 3488
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11422 3476 11428 3528
rect 11480 3516 11486 3528
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 11480 3488 11621 3516
rect 11480 3476 11486 3488
rect 11609 3485 11621 3488
rect 11655 3485 11667 3519
rect 11882 3516 11888 3528
rect 11795 3488 11888 3516
rect 11609 3479 11667 3485
rect 11882 3476 11888 3488
rect 11940 3516 11946 3528
rect 12158 3516 12164 3528
rect 11940 3488 12164 3516
rect 11940 3476 11946 3488
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 12250 3476 12256 3528
rect 12308 3516 12314 3528
rect 12437 3519 12495 3525
rect 12437 3516 12449 3519
rect 12308 3488 12449 3516
rect 12308 3476 12314 3488
rect 12437 3485 12449 3488
rect 12483 3485 12495 3519
rect 12710 3516 12716 3528
rect 12671 3488 12716 3516
rect 12437 3479 12495 3485
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 13403 3488 13860 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 10778 3448 10784 3460
rect 10739 3420 10784 3448
rect 10778 3408 10784 3420
rect 10836 3408 10842 3460
rect 10870 3408 10876 3460
rect 10928 3448 10934 3460
rect 10981 3451 11039 3457
rect 10981 3448 10993 3451
rect 10928 3420 10993 3448
rect 10928 3408 10934 3420
rect 10981 3417 10993 3420
rect 11027 3417 11039 3451
rect 10981 3411 11039 3417
rect 11072 3420 11376 3448
rect 11072 3380 11100 3420
rect 10612 3352 11100 3380
rect 10321 3343 10379 3349
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 11348 3380 11376 3420
rect 11514 3408 11520 3460
rect 11572 3448 11578 3460
rect 11974 3448 11980 3460
rect 11572 3420 11980 3448
rect 11572 3408 11578 3420
rect 11974 3408 11980 3420
rect 12032 3408 12038 3460
rect 13170 3408 13176 3460
rect 13228 3448 13234 3460
rect 13722 3448 13728 3460
rect 13228 3420 13728 3448
rect 13228 3408 13234 3420
rect 13722 3408 13728 3420
rect 13780 3408 13786 3460
rect 12535 3383 12593 3389
rect 12535 3380 12547 3383
rect 11204 3352 11249 3380
rect 11348 3352 12547 3380
rect 11204 3340 11210 3352
rect 12535 3349 12547 3352
rect 12581 3349 12593 3383
rect 12535 3343 12593 3349
rect 12621 3383 12679 3389
rect 12621 3349 12633 3383
rect 12667 3380 12679 3383
rect 13630 3380 13636 3392
rect 12667 3352 13636 3380
rect 12667 3349 12679 3352
rect 12621 3343 12679 3349
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 13832 3380 13860 3488
rect 13906 3476 13912 3528
rect 13964 3516 13970 3528
rect 14829 3519 14887 3525
rect 14829 3516 14841 3519
rect 13964 3488 14841 3516
rect 13964 3476 13970 3488
rect 14829 3485 14841 3488
rect 14875 3485 14887 3519
rect 14829 3479 14887 3485
rect 15657 3519 15715 3525
rect 15657 3485 15669 3519
rect 15703 3516 15715 3519
rect 16114 3516 16120 3528
rect 15703 3488 16120 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 14185 3451 14243 3457
rect 14185 3417 14197 3451
rect 14231 3448 14243 3451
rect 14458 3448 14464 3460
rect 14231 3420 14464 3448
rect 14231 3417 14243 3420
rect 14185 3411 14243 3417
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 16298 3380 16304 3392
rect 13832 3352 16304 3380
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 1104 3290 16836 3312
rect 1104 3238 4898 3290
rect 4950 3238 4962 3290
rect 5014 3238 5026 3290
rect 5078 3238 5090 3290
rect 5142 3238 5154 3290
rect 5206 3238 8846 3290
rect 8898 3238 8910 3290
rect 8962 3238 8974 3290
rect 9026 3238 9038 3290
rect 9090 3238 9102 3290
rect 9154 3238 12794 3290
rect 12846 3238 12858 3290
rect 12910 3238 12922 3290
rect 12974 3238 12986 3290
rect 13038 3238 13050 3290
rect 13102 3238 16836 3290
rect 1104 3216 16836 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3145 1639 3179
rect 1581 3139 1639 3145
rect 1596 3108 1624 3139
rect 2130 3136 2136 3188
rect 2188 3176 2194 3188
rect 2498 3176 2504 3188
rect 2188 3148 2504 3176
rect 2188 3136 2194 3148
rect 2498 3136 2504 3148
rect 2556 3176 2562 3188
rect 4614 3176 4620 3188
rect 2556 3148 4620 3176
rect 2556 3136 2562 3148
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 7006 3176 7012 3188
rect 6528 3148 7012 3176
rect 4700 3111 4758 3117
rect 1596 3080 2544 3108
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2516 3040 2544 3080
rect 2746 3080 4476 3108
rect 2590 3040 2596 3052
rect 2503 3012 2596 3040
rect 2590 3000 2596 3012
rect 2648 3040 2654 3052
rect 2746 3040 2774 3080
rect 4448 3052 4476 3080
rect 4700 3077 4712 3111
rect 4746 3108 4758 3111
rect 5442 3108 5448 3120
rect 4746 3080 5448 3108
rect 4746 3077 4758 3080
rect 4700 3071 4758 3077
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 2866 3049 2872 3052
rect 2860 3040 2872 3049
rect 2648 3012 2774 3040
rect 2827 3012 2872 3040
rect 2648 3000 2654 3012
rect 2860 3003 2872 3012
rect 2866 3000 2872 3003
rect 2924 3000 2930 3052
rect 4430 3040 4436 3052
rect 4391 3012 4436 3040
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 6528 3049 6556 3148
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 9766 3176 9772 3188
rect 7156 3148 9772 3176
rect 7156 3136 7162 3148
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10229 3179 10287 3185
rect 10229 3176 10241 3179
rect 10008 3148 10241 3176
rect 10008 3136 10014 3148
rect 10229 3145 10241 3148
rect 10275 3145 10287 3179
rect 10229 3139 10287 3145
rect 10502 3136 10508 3188
rect 10560 3176 10566 3188
rect 10870 3176 10876 3188
rect 10560 3148 10876 3176
rect 10560 3136 10566 3148
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11885 3179 11943 3185
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 12066 3176 12072 3188
rect 11931 3148 12072 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 12158 3136 12164 3188
rect 12216 3176 12222 3188
rect 12526 3176 12532 3188
rect 12216 3148 12532 3176
rect 12216 3136 12222 3148
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 13357 3179 13415 3185
rect 13357 3145 13369 3179
rect 13403 3176 13415 3179
rect 13722 3176 13728 3188
rect 13403 3148 13728 3176
rect 13403 3145 13415 3148
rect 13357 3139 13415 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 15289 3179 15347 3185
rect 15289 3176 15301 3179
rect 13872 3148 15301 3176
rect 13872 3136 13878 3148
rect 15289 3145 15301 3148
rect 15335 3145 15347 3179
rect 15289 3139 15347 3145
rect 15470 3136 15476 3188
rect 15528 3176 15534 3188
rect 16482 3176 16488 3188
rect 15528 3148 16488 3176
rect 15528 3136 15534 3148
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 6730 3108 6736 3120
rect 6691 3080 6736 3108
rect 6730 3068 6736 3080
rect 6788 3068 6794 3120
rect 7466 3068 7472 3120
rect 7524 3108 7530 3120
rect 8754 3108 8760 3120
rect 7524 3080 8760 3108
rect 7524 3068 7530 3080
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 9030 3068 9036 3120
rect 9088 3108 9094 3120
rect 9490 3108 9496 3120
rect 9088 3080 9496 3108
rect 9088 3068 9094 3080
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 9585 3111 9643 3117
rect 9585 3077 9597 3111
rect 9631 3108 9643 3111
rect 10042 3108 10048 3120
rect 9631 3080 10048 3108
rect 9631 3077 9643 3080
rect 9585 3071 9643 3077
rect 10042 3068 10048 3080
rect 10100 3068 10106 3120
rect 11514 3108 11520 3120
rect 11475 3080 11520 3108
rect 11514 3068 11520 3080
rect 11572 3068 11578 3120
rect 11701 3111 11759 3117
rect 11701 3077 11713 3111
rect 11747 3108 11759 3111
rect 12434 3108 12440 3120
rect 11747 3080 12440 3108
rect 11747 3077 11759 3080
rect 11701 3071 11759 3077
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 13538 3108 13544 3120
rect 12544 3080 13544 3108
rect 12544 3052 12572 3080
rect 13538 3068 13544 3080
rect 13596 3068 13602 3120
rect 13906 3108 13912 3120
rect 13867 3080 13912 3108
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 14090 3108 14096 3120
rect 14051 3080 14096 3108
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14476 3080 15516 3108
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6513 3043 6571 3049
rect 6513 3009 6525 3043
rect 6559 3009 6571 3043
rect 6513 3003 6571 3009
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 6871 3043 6929 3049
rect 6871 3009 6883 3043
rect 6917 3040 6929 3043
rect 6917 3012 7788 3040
rect 6917 3009 6929 3012
rect 6871 3003 6929 3009
rect 1486 2932 1492 2984
rect 1544 2972 1550 2984
rect 1765 2975 1823 2981
rect 1765 2972 1777 2975
rect 1544 2944 1777 2972
rect 1544 2932 1550 2944
rect 1765 2941 1777 2944
rect 1811 2941 1823 2975
rect 1765 2935 1823 2941
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2972 2099 2975
rect 2498 2972 2504 2984
rect 2087 2944 2504 2972
rect 2087 2941 2099 2944
rect 2041 2935 2099 2941
rect 1872 2836 1900 2935
rect 2498 2932 2504 2944
rect 2556 2932 2562 2984
rect 5442 2932 5448 2984
rect 5500 2972 5506 2984
rect 5718 2972 5724 2984
rect 5500 2944 5724 2972
rect 5500 2932 5506 2944
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 1946 2864 1952 2916
rect 2004 2904 2010 2916
rect 2130 2904 2136 2916
rect 2004 2876 2136 2904
rect 2004 2864 2010 2876
rect 2130 2864 2136 2876
rect 2188 2864 2194 2916
rect 3973 2907 4031 2913
rect 3973 2873 3985 2907
rect 4019 2904 4031 2907
rect 4154 2904 4160 2916
rect 4019 2876 4160 2904
rect 4019 2873 4031 2876
rect 3973 2867 4031 2873
rect 4154 2864 4160 2876
rect 4212 2864 4218 2916
rect 5534 2864 5540 2916
rect 5592 2904 5598 2916
rect 5813 2907 5871 2913
rect 5813 2904 5825 2907
rect 5592 2876 5825 2904
rect 5592 2864 5598 2876
rect 5813 2873 5825 2876
rect 5859 2873 5871 2907
rect 6380 2904 6408 3003
rect 6656 2972 6684 3003
rect 7558 2972 7564 2984
rect 6656 2944 7564 2972
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 7760 2972 7788 3012
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 7892 3012 7937 3040
rect 8588 3012 9720 3040
rect 7892 3000 7898 3012
rect 8588 2972 8616 3012
rect 7760 2944 8616 2972
rect 8662 2932 8668 2984
rect 8720 2972 8726 2984
rect 9306 2972 9312 2984
rect 8720 2944 9312 2972
rect 8720 2932 8726 2944
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 9692 2972 9720 3012
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 12345 3043 12403 3049
rect 12345 3040 12357 3043
rect 9824 3030 10088 3040
rect 10244 3030 12357 3040
rect 9824 3012 12357 3030
rect 9824 3000 9830 3012
rect 10060 3002 10272 3012
rect 12345 3009 12357 3012
rect 12391 3040 12403 3043
rect 12526 3040 12532 3052
rect 12391 3012 12532 3040
rect 12391 3009 12403 3012
rect 12345 3003 12403 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12621 3043 12679 3049
rect 12621 3009 12633 3043
rect 12667 3040 12679 3043
rect 12710 3040 12716 3052
rect 12667 3012 12716 3040
rect 12667 3009 12679 3012
rect 12621 3003 12679 3009
rect 12710 3000 12716 3012
rect 12768 3040 12774 3052
rect 13078 3040 13084 3052
rect 12768 3012 13084 3040
rect 12768 3000 12774 3012
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13262 3040 13268 3052
rect 13219 3012 13268 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3040 13507 3043
rect 13722 3040 13728 3052
rect 13495 3012 13728 3040
rect 13495 3009 13507 3012
rect 13449 3003 13507 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14185 3043 14243 3049
rect 14185 3009 14197 3043
rect 14231 3040 14243 3043
rect 14366 3040 14372 3052
rect 14231 3012 14372 3040
rect 14231 3009 14243 3012
rect 14185 3003 14243 3009
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 11054 2972 11060 2984
rect 9692 2944 11060 2972
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 13538 2932 13544 2984
rect 13596 2972 13602 2984
rect 14476 2972 14504 3080
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 14645 3043 14703 3049
rect 14645 3040 14657 3043
rect 14608 3012 14657 3040
rect 14608 3000 14614 3012
rect 14645 3009 14657 3012
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3040 14887 3043
rect 15378 3040 15384 3052
rect 14875 3012 15384 3040
rect 14875 3009 14887 3012
rect 14829 3003 14887 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 15488 3049 15516 3080
rect 15473 3043 15531 3049
rect 15473 3009 15485 3043
rect 15519 3009 15531 3043
rect 15473 3003 15531 3009
rect 15838 3000 15844 3052
rect 15896 3040 15902 3052
rect 15933 3043 15991 3049
rect 15933 3040 15945 3043
rect 15896 3012 15945 3040
rect 15896 3000 15902 3012
rect 15933 3009 15945 3012
rect 15979 3009 15991 3043
rect 15933 3003 15991 3009
rect 13596 2944 14504 2972
rect 13596 2932 13602 2944
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 14792 2944 16160 2972
rect 14792 2932 14798 2944
rect 8018 2904 8024 2916
rect 6380 2876 8024 2904
rect 5813 2867 5871 2873
rect 8018 2864 8024 2876
rect 8076 2864 8082 2916
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 12437 2907 12495 2913
rect 12437 2904 12449 2907
rect 9732 2876 12449 2904
rect 9732 2864 9738 2876
rect 12437 2873 12449 2876
rect 12483 2873 12495 2907
rect 12437 2867 12495 2873
rect 12802 2864 12808 2916
rect 12860 2904 12866 2916
rect 13173 2907 13231 2913
rect 13173 2904 13185 2907
rect 12860 2876 13185 2904
rect 12860 2864 12866 2876
rect 13173 2873 13185 2876
rect 13219 2904 13231 2907
rect 15102 2904 15108 2916
rect 13219 2876 15108 2904
rect 13219 2873 13231 2876
rect 13173 2867 13231 2873
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 16132 2913 16160 2944
rect 16117 2907 16175 2913
rect 16117 2873 16129 2907
rect 16163 2873 16175 2907
rect 16117 2867 16175 2873
rect 4062 2836 4068 2848
rect 1872 2808 4068 2836
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 7009 2839 7067 2845
rect 7009 2836 7021 2839
rect 5224 2808 7021 2836
rect 5224 2796 5230 2808
rect 7009 2805 7021 2808
rect 7055 2805 7067 2839
rect 7009 2799 7067 2805
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 10229 2839 10287 2845
rect 10229 2836 10241 2839
rect 8444 2808 10241 2836
rect 8444 2796 8450 2808
rect 10229 2805 10241 2808
rect 10275 2805 10287 2839
rect 10410 2836 10416 2848
rect 10371 2808 10416 2836
rect 10229 2799 10287 2805
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 10502 2796 10508 2848
rect 10560 2836 10566 2848
rect 10778 2836 10784 2848
rect 10560 2808 10784 2836
rect 10560 2796 10566 2808
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 11882 2836 11888 2848
rect 11296 2808 11888 2836
rect 11296 2796 11302 2808
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 12342 2796 12348 2848
rect 12400 2836 12406 2848
rect 13078 2836 13084 2848
rect 12400 2808 13084 2836
rect 12400 2796 12406 2808
rect 13078 2796 13084 2808
rect 13136 2836 13142 2848
rect 13722 2836 13728 2848
rect 13136 2808 13728 2836
rect 13136 2796 13142 2808
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 13814 2796 13820 2848
rect 13872 2836 13878 2848
rect 13909 2839 13967 2845
rect 13909 2836 13921 2839
rect 13872 2808 13921 2836
rect 13872 2796 13878 2808
rect 13909 2805 13921 2808
rect 13955 2805 13967 2839
rect 14642 2836 14648 2848
rect 14603 2808 14648 2836
rect 13909 2799 13967 2805
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 1104 2746 16836 2768
rect 1104 2694 2924 2746
rect 2976 2694 2988 2746
rect 3040 2694 3052 2746
rect 3104 2694 3116 2746
rect 3168 2694 3180 2746
rect 3232 2694 6872 2746
rect 6924 2694 6936 2746
rect 6988 2694 7000 2746
rect 7052 2694 7064 2746
rect 7116 2694 7128 2746
rect 7180 2694 10820 2746
rect 10872 2694 10884 2746
rect 10936 2694 10948 2746
rect 11000 2694 11012 2746
rect 11064 2694 11076 2746
rect 11128 2694 14768 2746
rect 14820 2694 14832 2746
rect 14884 2694 14896 2746
rect 14948 2694 14960 2746
rect 15012 2694 15024 2746
rect 15076 2694 16836 2746
rect 1104 2672 16836 2694
rect 2774 2632 2780 2644
rect 1412 2604 2780 2632
rect 1412 2505 1440 2604
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 3142 2592 3148 2644
rect 3200 2632 3206 2644
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 3200 2604 7573 2632
rect 3200 2592 3206 2604
rect 7561 2601 7573 2604
rect 7607 2632 7619 2635
rect 7834 2632 7840 2644
rect 7607 2604 7840 2632
rect 7607 2601 7619 2604
rect 7561 2595 7619 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8018 2632 8024 2644
rect 7979 2604 8024 2632
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 8202 2592 8208 2644
rect 8260 2632 8266 2644
rect 10134 2632 10140 2644
rect 8260 2604 10140 2632
rect 8260 2592 8266 2604
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 10744 2604 11713 2632
rect 10744 2592 10750 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 11701 2595 11759 2601
rect 11882 2592 11888 2644
rect 11940 2632 11946 2644
rect 11940 2604 13492 2632
rect 11940 2592 11946 2604
rect 2130 2524 2136 2576
rect 2188 2564 2194 2576
rect 3789 2567 3847 2573
rect 3789 2564 3801 2567
rect 2188 2536 3801 2564
rect 2188 2524 2194 2536
rect 3789 2533 3801 2536
rect 3835 2533 3847 2567
rect 3789 2527 3847 2533
rect 4062 2524 4068 2576
rect 4120 2564 4126 2576
rect 4120 2536 4568 2564
rect 4120 2524 4126 2536
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 1762 2496 1768 2508
rect 1719 2468 1768 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 1762 2456 1768 2468
rect 1820 2456 1826 2508
rect 2682 2456 2688 2508
rect 2740 2496 2746 2508
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 2740 2468 2789 2496
rect 2740 2456 2746 2468
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 2777 2459 2835 2465
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2465 4491 2499
rect 4540 2496 4568 2536
rect 5902 2524 5908 2576
rect 5960 2564 5966 2576
rect 8294 2564 8300 2576
rect 5960 2536 8300 2564
rect 5960 2524 5966 2536
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 8846 2524 8852 2576
rect 8904 2564 8910 2576
rect 11054 2564 11060 2576
rect 8904 2536 11060 2564
rect 8904 2524 8910 2536
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 11974 2564 11980 2576
rect 11195 2536 11980 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 11974 2524 11980 2536
rect 12032 2524 12038 2576
rect 12526 2524 12532 2576
rect 12584 2564 12590 2576
rect 13357 2567 13415 2573
rect 13357 2564 13369 2567
rect 12584 2536 13369 2564
rect 12584 2524 12590 2536
rect 13357 2533 13369 2536
rect 13403 2533 13415 2567
rect 13464 2564 13492 2604
rect 14182 2592 14188 2644
rect 14240 2632 14246 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 14240 2604 14289 2632
rect 14240 2592 14246 2604
rect 14277 2601 14289 2604
rect 14323 2601 14335 2635
rect 15562 2632 15568 2644
rect 14277 2595 14335 2601
rect 14384 2604 15568 2632
rect 14384 2564 14412 2604
rect 15562 2592 15568 2604
rect 15620 2592 15626 2644
rect 15841 2635 15899 2641
rect 15841 2601 15853 2635
rect 15887 2632 15899 2635
rect 16206 2632 16212 2644
rect 15887 2604 16212 2632
rect 15887 2601 15899 2604
rect 15841 2595 15899 2601
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 13464 2536 14412 2564
rect 13357 2527 13415 2533
rect 14918 2524 14924 2576
rect 14976 2564 14982 2576
rect 16482 2564 16488 2576
rect 14976 2536 16488 2564
rect 14976 2524 14982 2536
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 6178 2496 6184 2508
rect 4540 2468 6184 2496
rect 4433 2459 4491 2465
rect 1780 2360 1808 2456
rect 2866 2428 2872 2440
rect 2827 2400 2872 2428
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 4448 2428 4476 2459
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2496 7067 2499
rect 12066 2496 12072 2508
rect 7055 2468 11652 2496
rect 7055 2465 7067 2468
rect 7009 2459 7067 2465
rect 11624 2440 11652 2468
rect 11732 2468 12072 2496
rect 5626 2428 5632 2440
rect 4448 2400 5632 2428
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 6638 2428 6644 2440
rect 5776 2400 6644 2428
rect 5776 2388 5782 2400
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 7616 2400 7757 2428
rect 7616 2388 7622 2400
rect 7745 2397 7757 2400
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 8662 2388 8668 2440
rect 8720 2428 8726 2440
rect 9030 2428 9036 2440
rect 8720 2400 9036 2428
rect 8720 2388 8726 2400
rect 9030 2388 9036 2400
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 9401 2431 9459 2437
rect 9401 2428 9413 2431
rect 9272 2400 9413 2428
rect 9272 2388 9278 2400
rect 9401 2397 9413 2400
rect 9447 2397 9459 2431
rect 9401 2391 9459 2397
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 10045 2431 10103 2437
rect 10045 2428 10057 2431
rect 9916 2400 10057 2428
rect 9916 2388 9922 2400
rect 10045 2397 10057 2400
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2428 10379 2431
rect 10367 2400 10732 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 4249 2363 4307 2369
rect 4249 2360 4261 2363
rect 1780 2332 4261 2360
rect 4249 2329 4261 2332
rect 4295 2329 4307 2363
rect 4249 2323 4307 2329
rect 5261 2363 5319 2369
rect 5261 2329 5273 2363
rect 5307 2360 5319 2363
rect 10594 2360 10600 2372
rect 5307 2332 10600 2360
rect 5307 2329 5319 2332
rect 5261 2323 5319 2329
rect 10594 2320 10600 2332
rect 10652 2320 10658 2372
rect 10704 2360 10732 2400
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 10965 2431 11023 2437
rect 10836 2400 10881 2428
rect 10836 2388 10842 2400
rect 10965 2397 10977 2431
rect 11011 2397 11023 2431
rect 11606 2428 11612 2440
rect 11519 2400 11612 2428
rect 10965 2391 11023 2397
rect 10980 2360 11008 2391
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 11732 2360 11760 2468
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 12434 2496 12440 2508
rect 12216 2468 12440 2496
rect 12216 2456 12222 2468
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 12618 2496 12624 2508
rect 12544 2468 12624 2496
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 12544 2437 12572 2468
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 12805 2499 12863 2505
rect 12805 2465 12817 2499
rect 12851 2496 12863 2499
rect 16574 2496 16580 2508
rect 12851 2468 16580 2496
rect 12851 2465 12863 2468
rect 12805 2459 12863 2465
rect 16574 2456 16580 2468
rect 16632 2456 16638 2508
rect 12529 2431 12587 2437
rect 11848 2400 11893 2428
rect 11848 2388 11854 2400
rect 12529 2397 12541 2431
rect 12575 2397 12587 2431
rect 12710 2428 12716 2440
rect 12671 2400 12716 2428
rect 12529 2391 12587 2397
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 12986 2388 12992 2440
rect 13044 2388 13050 2440
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 13136 2400 13277 2428
rect 13136 2388 13142 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 13630 2428 13636 2440
rect 13587 2400 13636 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 14182 2428 14188 2440
rect 14143 2400 14188 2428
rect 14182 2388 14188 2400
rect 14240 2428 14246 2440
rect 14918 2428 14924 2440
rect 14240 2400 14924 2428
rect 14240 2388 14246 2400
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 15194 2428 15200 2440
rect 15059 2400 15200 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 15746 2388 15752 2440
rect 15804 2428 15810 2440
rect 15841 2431 15899 2437
rect 15841 2428 15853 2431
rect 15804 2400 15853 2428
rect 15804 2388 15810 2400
rect 15841 2397 15853 2400
rect 15887 2397 15899 2431
rect 16022 2428 16028 2440
rect 15983 2400 16028 2428
rect 15841 2391 15899 2397
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 13004 2360 13032 2388
rect 10704 2332 10916 2360
rect 10980 2332 11760 2360
rect 11799 2332 13032 2360
rect 13449 2363 13507 2369
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 3970 2292 3976 2304
rect 3283 2264 3976 2292
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 4157 2295 4215 2301
rect 4157 2261 4169 2295
rect 4203 2292 4215 2295
rect 4430 2292 4436 2304
rect 4203 2264 4436 2292
rect 4203 2261 4215 2264
rect 4157 2255 4215 2261
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 4614 2252 4620 2304
rect 4672 2292 4678 2304
rect 8846 2292 8852 2304
rect 4672 2264 8852 2292
rect 4672 2252 4678 2264
rect 8846 2252 8852 2264
rect 8904 2252 8910 2304
rect 8941 2295 8999 2301
rect 8941 2261 8953 2295
rect 8987 2292 8999 2295
rect 9214 2292 9220 2304
rect 8987 2264 9220 2292
rect 8987 2261 8999 2264
rect 8941 2255 8999 2261
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 9309 2295 9367 2301
rect 9309 2261 9321 2295
rect 9355 2292 9367 2295
rect 9490 2292 9496 2304
rect 9355 2264 9496 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 9490 2252 9496 2264
rect 9548 2252 9554 2304
rect 9861 2295 9919 2301
rect 9861 2261 9873 2295
rect 9907 2292 9919 2295
rect 10042 2292 10048 2304
rect 9907 2264 10048 2292
rect 9907 2261 9919 2264
rect 9861 2255 9919 2261
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10226 2252 10232 2304
rect 10284 2292 10290 2304
rect 10888 2292 10916 2332
rect 10962 2292 10968 2304
rect 10284 2264 10329 2292
rect 10888 2264 10968 2292
rect 10284 2252 10290 2264
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11054 2252 11060 2304
rect 11112 2292 11118 2304
rect 11799 2292 11827 2332
rect 13449 2329 13461 2363
rect 13495 2329 13507 2363
rect 13449 2323 13507 2329
rect 11112 2264 11827 2292
rect 11112 2252 11118 2264
rect 12434 2252 12440 2304
rect 12492 2292 12498 2304
rect 12802 2292 12808 2304
rect 12492 2264 12808 2292
rect 12492 2252 12498 2264
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13464 2292 13492 2323
rect 14826 2292 14832 2304
rect 12952 2264 13492 2292
rect 14787 2264 14832 2292
rect 12952 2252 12958 2264
rect 14826 2252 14832 2264
rect 14884 2252 14890 2304
rect 1104 2202 16836 2224
rect 1104 2150 4898 2202
rect 4950 2150 4962 2202
rect 5014 2150 5026 2202
rect 5078 2150 5090 2202
rect 5142 2150 5154 2202
rect 5206 2150 8846 2202
rect 8898 2150 8910 2202
rect 8962 2150 8974 2202
rect 9026 2150 9038 2202
rect 9090 2150 9102 2202
rect 9154 2150 12794 2202
rect 12846 2150 12858 2202
rect 12910 2150 12922 2202
rect 12974 2150 12986 2202
rect 13038 2150 13050 2202
rect 13102 2150 16836 2202
rect 1104 2128 16836 2150
rect 3053 2091 3111 2097
rect 3053 2057 3065 2091
rect 3099 2088 3111 2091
rect 3789 2091 3847 2097
rect 3789 2088 3801 2091
rect 3099 2060 3801 2088
rect 3099 2057 3111 2060
rect 3053 2051 3111 2057
rect 3789 2057 3801 2060
rect 3835 2057 3847 2091
rect 5813 2091 5871 2097
rect 3789 2051 3847 2057
rect 3896 2060 5672 2088
rect 1026 1980 1032 2032
rect 1084 2020 1090 2032
rect 1084 1992 2176 2020
rect 1084 1980 1090 1992
rect 2041 1955 2099 1961
rect 2041 1921 2053 1955
rect 2087 1952 2099 1955
rect 2148 1952 2176 1992
rect 3418 1980 3424 2032
rect 3476 2020 3482 2032
rect 3896 2020 3924 2060
rect 4154 2020 4160 2032
rect 3476 1992 3924 2020
rect 4115 1992 4160 2020
rect 3476 1980 3482 1992
rect 4154 1980 4160 1992
rect 4212 1980 4218 2032
rect 4798 1980 4804 2032
rect 4856 2020 4862 2032
rect 5445 2023 5503 2029
rect 5445 2020 5457 2023
rect 4856 1992 5457 2020
rect 4856 1980 4862 1992
rect 5445 1989 5457 1992
rect 5491 1989 5503 2023
rect 5445 1983 5503 1989
rect 2222 1952 2228 1964
rect 2087 1924 2228 1952
rect 2087 1921 2099 1924
rect 2041 1915 2099 1921
rect 2222 1912 2228 1924
rect 2280 1912 2286 1964
rect 4246 1952 4252 1964
rect 4159 1924 4252 1952
rect 4246 1912 4252 1924
rect 4304 1952 4310 1964
rect 5166 1952 5172 1964
rect 4304 1924 5172 1952
rect 4304 1912 4310 1924
rect 5166 1912 5172 1924
rect 5224 1912 5230 1964
rect 5261 1955 5319 1961
rect 5261 1921 5273 1955
rect 5307 1921 5319 1955
rect 5534 1952 5540 1964
rect 5495 1924 5540 1952
rect 5261 1915 5319 1921
rect 1857 1887 1915 1893
rect 1857 1853 1869 1887
rect 1903 1853 1915 1887
rect 1857 1847 1915 1853
rect 1872 1816 1900 1847
rect 1946 1844 1952 1896
rect 2004 1884 2010 1896
rect 2133 1887 2191 1893
rect 2004 1856 2049 1884
rect 2004 1844 2010 1856
rect 2133 1853 2145 1887
rect 2179 1884 2191 1887
rect 2682 1884 2688 1896
rect 2179 1856 2688 1884
rect 2179 1853 2191 1856
rect 2133 1847 2191 1853
rect 2682 1844 2688 1856
rect 2740 1844 2746 1896
rect 4062 1884 4068 1896
rect 3160 1856 4068 1884
rect 3160 1816 3188 1856
rect 4062 1844 4068 1856
rect 4120 1884 4126 1896
rect 4433 1887 4491 1893
rect 4433 1884 4445 1887
rect 4120 1856 4445 1884
rect 4120 1844 4126 1856
rect 4433 1853 4445 1856
rect 4479 1884 4491 1887
rect 5074 1884 5080 1896
rect 4479 1856 5080 1884
rect 4479 1853 4491 1856
rect 4433 1847 4491 1853
rect 5074 1844 5080 1856
rect 5132 1844 5138 1896
rect 5276 1884 5304 1915
rect 5534 1912 5540 1924
rect 5592 1912 5598 1964
rect 5644 1961 5672 2060
rect 5813 2057 5825 2091
rect 5859 2088 5871 2091
rect 5994 2088 6000 2100
rect 5859 2060 6000 2088
rect 5859 2057 5871 2060
rect 5813 2051 5871 2057
rect 5994 2048 6000 2060
rect 6052 2048 6058 2100
rect 9766 2088 9772 2100
rect 6196 2060 9772 2088
rect 5629 1955 5687 1961
rect 5629 1921 5641 1955
rect 5675 1921 5687 1955
rect 5629 1915 5687 1921
rect 6196 1884 6224 2060
rect 9766 2048 9772 2060
rect 9824 2048 9830 2100
rect 10042 2048 10048 2100
rect 10100 2088 10106 2100
rect 11882 2088 11888 2100
rect 10100 2060 10180 2088
rect 10100 2048 10106 2060
rect 6270 1980 6276 2032
rect 6328 2020 6334 2032
rect 6365 2023 6423 2029
rect 6365 2020 6377 2023
rect 6328 1992 6377 2020
rect 6328 1980 6334 1992
rect 6365 1989 6377 1992
rect 6411 1989 6423 2023
rect 7006 2020 7012 2032
rect 6365 1983 6423 1989
rect 6564 1992 7012 2020
rect 6564 1961 6592 1992
rect 7006 1980 7012 1992
rect 7064 1980 7070 2032
rect 8570 2020 8576 2032
rect 7116 1992 8576 2020
rect 6549 1955 6607 1961
rect 6549 1952 6561 1955
rect 5276 1856 6224 1884
rect 6472 1924 6561 1952
rect 1872 1788 3188 1816
rect 3237 1819 3295 1825
rect 3237 1785 3249 1819
rect 3283 1816 3295 1819
rect 3786 1816 3792 1828
rect 3283 1788 3792 1816
rect 3283 1785 3295 1788
rect 3237 1779 3295 1785
rect 3786 1776 3792 1788
rect 3844 1776 3850 1828
rect 4246 1776 4252 1828
rect 4304 1816 4310 1828
rect 6472 1816 6500 1924
rect 6549 1921 6561 1924
rect 6595 1921 6607 1955
rect 6549 1915 6607 1921
rect 6641 1955 6699 1961
rect 6641 1921 6653 1955
rect 6687 1952 6699 1955
rect 6730 1952 6736 1964
rect 6687 1924 6736 1952
rect 6687 1921 6699 1924
rect 6641 1915 6699 1921
rect 6730 1912 6736 1924
rect 6788 1912 6794 1964
rect 7116 1961 7144 1992
rect 8570 1980 8576 1992
rect 8628 1980 8634 2032
rect 9030 1980 9036 2032
rect 9088 2020 9094 2032
rect 9088 1992 10088 2020
rect 9088 1980 9094 1992
rect 7101 1955 7159 1961
rect 7101 1921 7113 1955
rect 7147 1921 7159 1955
rect 7101 1915 7159 1921
rect 7368 1955 7426 1961
rect 7368 1921 7380 1955
rect 7414 1952 7426 1955
rect 8941 1955 8999 1961
rect 7414 1924 8892 1952
rect 7414 1921 7426 1924
rect 7368 1915 7426 1921
rect 8864 1884 8892 1924
rect 8941 1921 8953 1955
rect 8987 1952 8999 1955
rect 9674 1952 9680 1964
rect 8987 1924 9680 1952
rect 8987 1921 8999 1924
rect 8941 1915 8999 1921
rect 9674 1912 9680 1924
rect 9732 1912 9738 1964
rect 9858 1952 9864 1964
rect 9819 1924 9864 1952
rect 9858 1912 9864 1924
rect 9916 1912 9922 1964
rect 10060 1961 10088 1992
rect 10045 1955 10103 1961
rect 10045 1921 10057 1955
rect 10091 1921 10103 1955
rect 10152 1952 10180 2060
rect 10428 2060 11888 2088
rect 10226 1980 10232 2032
rect 10284 2020 10290 2032
rect 10284 1992 10329 2020
rect 10284 1980 10290 1992
rect 10321 1955 10379 1961
rect 10321 1952 10333 1955
rect 10152 1924 10333 1952
rect 10045 1915 10103 1921
rect 10321 1921 10333 1924
rect 10367 1921 10379 1955
rect 10321 1915 10379 1921
rect 8864 1856 9536 1884
rect 7098 1816 7104 1828
rect 4304 1788 6500 1816
rect 6528 1788 7104 1816
rect 4304 1776 4310 1788
rect 1673 1751 1731 1757
rect 1673 1717 1685 1751
rect 1719 1748 1731 1751
rect 2774 1748 2780 1760
rect 1719 1720 2780 1748
rect 1719 1717 1731 1720
rect 1673 1711 1731 1717
rect 2774 1708 2780 1720
rect 2832 1708 2838 1760
rect 3053 1751 3111 1757
rect 3053 1717 3065 1751
rect 3099 1748 3111 1751
rect 3326 1748 3332 1760
rect 3099 1720 3332 1748
rect 3099 1717 3111 1720
rect 3053 1711 3111 1717
rect 3326 1708 3332 1720
rect 3384 1748 3390 1760
rect 6528 1748 6556 1788
rect 7098 1776 7104 1788
rect 7156 1776 7162 1828
rect 8294 1776 8300 1828
rect 8352 1816 8358 1828
rect 8481 1819 8539 1825
rect 8481 1816 8493 1819
rect 8352 1788 8493 1816
rect 8352 1776 8358 1788
rect 8481 1785 8493 1788
rect 8527 1785 8539 1819
rect 8481 1779 8539 1785
rect 8570 1776 8576 1828
rect 8628 1816 8634 1828
rect 9508 1816 9536 1856
rect 9766 1844 9772 1896
rect 9824 1884 9830 1896
rect 10428 1884 10456 2060
rect 11882 2048 11888 2060
rect 11940 2048 11946 2100
rect 12066 2048 12072 2100
rect 12124 2088 12130 2100
rect 12713 2091 12771 2097
rect 12713 2088 12725 2091
rect 12124 2060 12725 2088
rect 12124 2048 12130 2060
rect 12713 2057 12725 2060
rect 12759 2088 12771 2091
rect 12759 2060 13492 2088
rect 12759 2057 12771 2060
rect 12713 2051 12771 2057
rect 10870 1980 10876 2032
rect 10928 2020 10934 2032
rect 10928 1992 10973 2020
rect 10928 1980 10934 1992
rect 11330 1980 11336 2032
rect 11388 2020 11394 2032
rect 12158 2020 12164 2032
rect 11388 1992 12164 2020
rect 11388 1980 11394 1992
rect 12158 1980 12164 1992
rect 12216 1980 12222 2032
rect 12802 1980 12808 2032
rect 12860 2020 12866 2032
rect 13262 2020 13268 2032
rect 12860 1992 13268 2020
rect 12860 1980 12866 1992
rect 13262 1980 13268 1992
rect 13320 2020 13326 2032
rect 13320 1992 13400 2020
rect 13320 1980 13326 1992
rect 10778 1952 10784 1964
rect 10739 1924 10784 1952
rect 10778 1912 10784 1924
rect 10836 1912 10842 1964
rect 10965 1955 11023 1961
rect 10965 1921 10977 1955
rect 11011 1921 11023 1955
rect 10965 1915 11023 1921
rect 9824 1856 10456 1884
rect 9824 1844 9830 1856
rect 10686 1844 10692 1896
rect 10744 1884 10750 1896
rect 10980 1884 11008 1915
rect 11146 1912 11152 1964
rect 11204 1952 11210 1964
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 11204 1924 11529 1952
rect 11204 1912 11210 1924
rect 11517 1921 11529 1924
rect 11563 1921 11575 1955
rect 11517 1915 11575 1921
rect 11701 1955 11759 1961
rect 11701 1921 11713 1955
rect 11747 1921 11759 1955
rect 11882 1952 11888 1964
rect 11843 1924 11888 1952
rect 11701 1915 11759 1921
rect 10744 1856 11008 1884
rect 10744 1844 10750 1856
rect 11330 1844 11336 1896
rect 11388 1884 11394 1896
rect 11716 1884 11744 1915
rect 11882 1912 11888 1924
rect 11940 1912 11946 1964
rect 12342 1952 12348 1964
rect 12303 1924 12348 1952
rect 12342 1912 12348 1924
rect 12400 1912 12406 1964
rect 12434 1912 12440 1964
rect 12492 1952 12498 1964
rect 12492 1924 12537 1952
rect 12492 1912 12498 1924
rect 12618 1912 12624 1964
rect 12676 1952 12682 1964
rect 13372 1961 13400 1992
rect 13173 1955 13231 1961
rect 13173 1952 13185 1955
rect 12676 1924 13185 1952
rect 12676 1912 12682 1924
rect 13173 1921 13185 1924
rect 13219 1921 13231 1955
rect 13173 1915 13231 1921
rect 13357 1955 13415 1961
rect 13357 1921 13369 1955
rect 13403 1921 13415 1955
rect 13464 1952 13492 2060
rect 13722 2048 13728 2100
rect 13780 2088 13786 2100
rect 14921 2091 14979 2097
rect 14921 2088 14933 2091
rect 13780 2060 14933 2088
rect 13780 2048 13786 2060
rect 14921 2057 14933 2060
rect 14967 2057 14979 2091
rect 14921 2051 14979 2057
rect 15470 2048 15476 2100
rect 15528 2088 15534 2100
rect 15565 2091 15623 2097
rect 15565 2088 15577 2091
rect 15528 2060 15577 2088
rect 15528 2048 15534 2060
rect 15565 2057 15577 2060
rect 15611 2057 15623 2091
rect 15565 2051 15623 2057
rect 13998 1980 14004 2032
rect 14056 2020 14062 2032
rect 14217 2023 14275 2029
rect 14056 1992 14101 2020
rect 14056 1980 14062 1992
rect 14217 1989 14229 2023
rect 14263 2020 14275 2023
rect 14458 2020 14464 2032
rect 14263 1992 14464 2020
rect 14263 1989 14275 1992
rect 14217 1983 14275 1989
rect 14458 1980 14464 1992
rect 14516 1980 14522 2032
rect 14829 1955 14887 1961
rect 14829 1952 14841 1955
rect 13464 1924 14841 1952
rect 13357 1915 13415 1921
rect 14829 1921 14841 1924
rect 14875 1921 14887 1955
rect 15010 1952 15016 1964
rect 14971 1924 15016 1952
rect 14829 1915 14887 1921
rect 15010 1912 15016 1924
rect 15068 1912 15074 1964
rect 15473 1955 15531 1961
rect 15473 1921 15485 1955
rect 15519 1921 15531 1955
rect 15473 1915 15531 1921
rect 11388 1856 11744 1884
rect 11388 1844 11394 1856
rect 10502 1816 10508 1828
rect 8628 1788 9444 1816
rect 9508 1788 10508 1816
rect 8628 1776 8634 1788
rect 3384 1720 6556 1748
rect 6641 1751 6699 1757
rect 3384 1708 3390 1720
rect 6641 1717 6653 1751
rect 6687 1748 6699 1751
rect 9122 1748 9128 1760
rect 6687 1720 9128 1748
rect 6687 1717 6699 1720
rect 6641 1711 6699 1717
rect 9122 1708 9128 1720
rect 9180 1708 9186 1760
rect 9217 1751 9275 1757
rect 9217 1717 9229 1751
rect 9263 1748 9275 1751
rect 9306 1748 9312 1760
rect 9263 1720 9312 1748
rect 9263 1717 9275 1720
rect 9217 1711 9275 1717
rect 9306 1708 9312 1720
rect 9364 1708 9370 1760
rect 9416 1757 9444 1788
rect 10502 1776 10508 1788
rect 10560 1776 10566 1828
rect 11716 1816 11744 1856
rect 11790 1844 11796 1896
rect 11848 1884 11854 1896
rect 13078 1884 13084 1896
rect 11848 1856 13084 1884
rect 11848 1844 11854 1856
rect 13078 1844 13084 1856
rect 13136 1844 13142 1896
rect 14090 1844 14096 1896
rect 14148 1884 14154 1896
rect 15488 1884 15516 1915
rect 14148 1856 15516 1884
rect 14148 1844 14154 1856
rect 12066 1816 12072 1828
rect 11716 1788 12072 1816
rect 12066 1776 12072 1788
rect 12124 1776 12130 1828
rect 12158 1776 12164 1828
rect 12216 1816 12222 1828
rect 13265 1819 13323 1825
rect 13265 1816 13277 1819
rect 12216 1788 13277 1816
rect 12216 1776 12222 1788
rect 13265 1785 13277 1788
rect 13311 1785 13323 1819
rect 13265 1779 13323 1785
rect 13446 1776 13452 1828
rect 13504 1816 13510 1828
rect 13722 1816 13728 1828
rect 13504 1788 13728 1816
rect 13504 1776 13510 1788
rect 13722 1776 13728 1788
rect 13780 1776 13786 1828
rect 9401 1751 9459 1757
rect 9401 1717 9413 1751
rect 9447 1748 9459 1751
rect 10962 1748 10968 1760
rect 9447 1720 10968 1748
rect 9447 1717 9459 1720
rect 9401 1711 9459 1717
rect 10962 1708 10968 1720
rect 11020 1708 11026 1760
rect 12529 1751 12587 1757
rect 12529 1717 12541 1751
rect 12575 1748 12587 1751
rect 12986 1748 12992 1760
rect 12575 1720 12992 1748
rect 12575 1717 12587 1720
rect 12529 1711 12587 1717
rect 12986 1708 12992 1720
rect 13044 1708 13050 1760
rect 13538 1708 13544 1760
rect 13596 1748 13602 1760
rect 14185 1751 14243 1757
rect 14185 1748 14197 1751
rect 13596 1720 14197 1748
rect 13596 1708 13602 1720
rect 14185 1717 14197 1720
rect 14231 1717 14243 1751
rect 14185 1711 14243 1717
rect 14369 1751 14427 1757
rect 14369 1717 14381 1751
rect 14415 1748 14427 1751
rect 17310 1748 17316 1760
rect 14415 1720 17316 1748
rect 14415 1717 14427 1720
rect 14369 1711 14427 1717
rect 17310 1708 17316 1720
rect 17368 1708 17374 1760
rect 1104 1658 16836 1680
rect 1104 1606 2924 1658
rect 2976 1606 2988 1658
rect 3040 1606 3052 1658
rect 3104 1606 3116 1658
rect 3168 1606 3180 1658
rect 3232 1606 6872 1658
rect 6924 1606 6936 1658
rect 6988 1606 7000 1658
rect 7052 1606 7064 1658
rect 7116 1606 7128 1658
rect 7180 1606 10820 1658
rect 10872 1606 10884 1658
rect 10936 1606 10948 1658
rect 11000 1606 11012 1658
rect 11064 1606 11076 1658
rect 11128 1606 14768 1658
rect 14820 1606 14832 1658
rect 14884 1606 14896 1658
rect 14948 1606 14960 1658
rect 15012 1606 15024 1658
rect 15076 1606 16836 1658
rect 1104 1584 16836 1606
rect 1670 1504 1676 1556
rect 1728 1544 1734 1556
rect 1857 1547 1915 1553
rect 1857 1544 1869 1547
rect 1728 1516 1869 1544
rect 1728 1504 1734 1516
rect 1857 1513 1869 1516
rect 1903 1513 1915 1547
rect 1857 1507 1915 1513
rect 2777 1547 2835 1553
rect 2777 1513 2789 1547
rect 2823 1544 2835 1547
rect 4157 1547 4215 1553
rect 2823 1516 4108 1544
rect 2823 1513 2835 1516
rect 2777 1507 2835 1513
rect 3234 1476 3240 1488
rect 2746 1448 3240 1476
rect 2746 1408 2774 1448
rect 3234 1436 3240 1448
rect 3292 1436 3298 1488
rect 4080 1476 4108 1516
rect 4157 1513 4169 1547
rect 4203 1544 4215 1547
rect 4203 1516 5028 1544
rect 4203 1513 4215 1516
rect 4157 1507 4215 1513
rect 4522 1476 4528 1488
rect 4080 1448 4528 1476
rect 4522 1436 4528 1448
rect 4580 1436 4586 1488
rect 4706 1436 4712 1488
rect 4764 1476 4770 1488
rect 5000 1485 5028 1516
rect 5074 1504 5080 1556
rect 5132 1544 5138 1556
rect 6454 1544 6460 1556
rect 5132 1516 6460 1544
rect 5132 1504 5138 1516
rect 6454 1504 6460 1516
rect 6512 1504 6518 1556
rect 6549 1547 6607 1553
rect 6549 1513 6561 1547
rect 6595 1544 6607 1547
rect 6730 1544 6736 1556
rect 6595 1516 6736 1544
rect 6595 1513 6607 1516
rect 6549 1507 6607 1513
rect 6730 1504 6736 1516
rect 6788 1504 6794 1556
rect 8205 1547 8263 1553
rect 8205 1544 8217 1547
rect 6840 1516 8217 1544
rect 4893 1479 4951 1485
rect 4893 1476 4905 1479
rect 4764 1448 4905 1476
rect 4764 1436 4770 1448
rect 4893 1445 4905 1448
rect 4939 1445 4951 1479
rect 4893 1439 4951 1445
rect 4985 1479 5043 1485
rect 4985 1445 4997 1479
rect 5031 1476 5043 1479
rect 5442 1476 5448 1488
rect 5031 1448 5448 1476
rect 5031 1445 5043 1448
rect 4985 1439 5043 1445
rect 5442 1436 5448 1448
rect 5500 1436 5506 1488
rect 5629 1479 5687 1485
rect 5629 1445 5641 1479
rect 5675 1476 5687 1479
rect 6362 1476 6368 1488
rect 5675 1448 6368 1476
rect 5675 1445 5687 1448
rect 5629 1439 5687 1445
rect 6362 1436 6368 1448
rect 6420 1436 6426 1488
rect 6638 1436 6644 1488
rect 6696 1476 6702 1488
rect 6840 1476 6868 1516
rect 8205 1513 8217 1516
rect 8251 1513 8263 1547
rect 8205 1507 8263 1513
rect 8478 1504 8484 1556
rect 8536 1544 8542 1556
rect 8938 1544 8944 1556
rect 8536 1516 8944 1544
rect 8536 1504 8542 1516
rect 8938 1504 8944 1516
rect 8996 1504 9002 1556
rect 9490 1544 9496 1556
rect 9048 1516 9496 1544
rect 6696 1448 6868 1476
rect 7653 1479 7711 1485
rect 6696 1436 6702 1448
rect 7653 1445 7665 1479
rect 7699 1476 7711 1479
rect 9048 1476 9076 1516
rect 9490 1504 9496 1516
rect 9548 1504 9554 1556
rect 9950 1504 9956 1556
rect 10008 1544 10014 1556
rect 10045 1547 10103 1553
rect 10045 1544 10057 1547
rect 10008 1516 10057 1544
rect 10008 1504 10014 1516
rect 10045 1513 10057 1516
rect 10091 1513 10103 1547
rect 10045 1507 10103 1513
rect 10502 1504 10508 1556
rect 10560 1544 10566 1556
rect 11514 1544 11520 1556
rect 10560 1516 11520 1544
rect 10560 1504 10566 1516
rect 11514 1504 11520 1516
rect 11572 1504 11578 1556
rect 11698 1544 11704 1556
rect 11659 1516 11704 1544
rect 11698 1504 11704 1516
rect 11756 1504 11762 1556
rect 11790 1504 11796 1556
rect 11848 1544 11854 1556
rect 12066 1544 12072 1556
rect 11848 1516 12072 1544
rect 11848 1504 11854 1516
rect 12066 1504 12072 1516
rect 12124 1504 12130 1556
rect 13262 1544 13268 1556
rect 12360 1516 13124 1544
rect 13223 1516 13268 1544
rect 7699 1448 9076 1476
rect 7699 1445 7711 1448
rect 7653 1439 7711 1445
rect 9122 1436 9128 1488
rect 9180 1476 9186 1488
rect 12360 1476 12388 1516
rect 9180 1448 12388 1476
rect 12437 1479 12495 1485
rect 9180 1436 9186 1448
rect 12437 1445 12449 1479
rect 12483 1445 12495 1479
rect 12437 1439 12495 1445
rect 2700 1380 2774 1408
rect 3789 1411 3847 1417
rect 2038 1340 2044 1352
rect 1999 1312 2044 1340
rect 2038 1300 2044 1312
rect 2096 1300 2102 1352
rect 2225 1343 2283 1349
rect 2225 1309 2237 1343
rect 2271 1309 2283 1343
rect 2225 1303 2283 1309
rect 566 1232 572 1284
rect 624 1272 630 1284
rect 2240 1272 2268 1303
rect 2314 1300 2320 1352
rect 2372 1340 2378 1352
rect 2372 1312 2417 1340
rect 2372 1300 2378 1312
rect 624 1244 2268 1272
rect 624 1232 630 1244
rect 750 1164 756 1216
rect 808 1204 814 1216
rect 2700 1204 2728 1380
rect 3789 1377 3801 1411
rect 3835 1408 3847 1411
rect 4246 1408 4252 1420
rect 3835 1380 4252 1408
rect 3835 1377 3847 1380
rect 3789 1371 3847 1377
rect 4246 1368 4252 1380
rect 4304 1368 4310 1420
rect 4338 1368 4344 1420
rect 4396 1408 4402 1420
rect 12452 1408 12480 1439
rect 13096 1408 13124 1516
rect 13262 1504 13268 1516
rect 13320 1504 13326 1556
rect 14182 1504 14188 1556
rect 14240 1544 14246 1556
rect 14277 1547 14335 1553
rect 14277 1544 14289 1547
rect 14240 1516 14289 1544
rect 14240 1504 14246 1516
rect 14277 1513 14289 1516
rect 14323 1513 14335 1547
rect 14277 1507 14335 1513
rect 14458 1504 14464 1556
rect 14516 1544 14522 1556
rect 17402 1544 17408 1556
rect 14516 1516 17408 1544
rect 14516 1504 14522 1516
rect 17402 1504 17408 1516
rect 17460 1504 17466 1556
rect 13170 1436 13176 1488
rect 13228 1476 13234 1488
rect 15197 1479 15255 1485
rect 15197 1476 15209 1479
rect 13228 1448 15209 1476
rect 13228 1436 13234 1448
rect 15197 1445 15209 1448
rect 15243 1445 15255 1479
rect 15197 1439 15255 1445
rect 13630 1408 13636 1420
rect 4396 1380 12480 1408
rect 12550 1380 12756 1408
rect 13096 1380 13636 1408
rect 4396 1368 4402 1380
rect 2958 1340 2964 1352
rect 2919 1312 2964 1340
rect 2958 1300 2964 1312
rect 3016 1300 3022 1352
rect 3234 1340 3240 1352
rect 3195 1312 3240 1340
rect 3234 1300 3240 1312
rect 3292 1300 3298 1352
rect 3973 1343 4031 1349
rect 3973 1309 3985 1343
rect 4019 1340 4031 1343
rect 4062 1340 4068 1352
rect 4019 1312 4068 1340
rect 4019 1309 4031 1312
rect 3973 1303 4031 1309
rect 4062 1300 4068 1312
rect 4120 1300 4126 1352
rect 4801 1343 4859 1349
rect 4801 1309 4813 1343
rect 4847 1309 4859 1343
rect 4801 1303 4859 1309
rect 5077 1343 5135 1349
rect 5077 1309 5089 1343
rect 5123 1340 5135 1343
rect 5166 1340 5172 1352
rect 5123 1312 5172 1340
rect 5123 1309 5135 1312
rect 5077 1303 5135 1309
rect 3142 1204 3148 1216
rect 808 1176 2728 1204
rect 3103 1176 3148 1204
rect 808 1164 814 1176
rect 3142 1164 3148 1176
rect 3200 1164 3206 1216
rect 4614 1204 4620 1216
rect 4575 1176 4620 1204
rect 4614 1164 4620 1176
rect 4672 1164 4678 1216
rect 4816 1204 4844 1303
rect 5166 1300 5172 1312
rect 5224 1300 5230 1352
rect 5813 1343 5871 1349
rect 5813 1309 5825 1343
rect 5859 1340 5871 1343
rect 6638 1340 6644 1352
rect 5859 1312 6644 1340
rect 5859 1309 5871 1312
rect 5813 1303 5871 1309
rect 6638 1300 6644 1312
rect 6696 1300 6702 1352
rect 6822 1340 6828 1352
rect 6783 1312 6828 1340
rect 6822 1300 6828 1312
rect 6880 1300 6886 1352
rect 8386 1340 8392 1352
rect 8347 1312 8392 1340
rect 8386 1300 8392 1312
rect 8444 1300 8450 1352
rect 8478 1300 8484 1352
rect 8536 1340 8542 1352
rect 9030 1340 9036 1352
rect 8536 1312 9036 1340
rect 8536 1300 8542 1312
rect 9030 1300 9036 1312
rect 9088 1340 9094 1352
rect 9125 1343 9183 1349
rect 9125 1340 9137 1343
rect 9088 1312 9137 1340
rect 9088 1300 9094 1312
rect 9125 1309 9137 1312
rect 9171 1309 9183 1343
rect 9125 1303 9183 1309
rect 9401 1343 9459 1349
rect 9401 1309 9413 1343
rect 9447 1340 9459 1343
rect 10781 1343 10839 1349
rect 9447 1312 10640 1340
rect 9447 1309 9459 1312
rect 9401 1303 9459 1309
rect 5994 1232 6000 1284
rect 6052 1272 6058 1284
rect 6365 1275 6423 1281
rect 6365 1272 6377 1275
rect 6052 1244 6377 1272
rect 6052 1232 6058 1244
rect 6365 1241 6377 1244
rect 6411 1241 6423 1275
rect 6546 1272 6552 1284
rect 6507 1244 6552 1272
rect 6365 1235 6423 1241
rect 6546 1232 6552 1244
rect 6604 1232 6610 1284
rect 7285 1275 7343 1281
rect 7285 1241 7297 1275
rect 7331 1272 7343 1275
rect 8662 1272 8668 1284
rect 7331 1244 8668 1272
rect 7331 1241 7343 1244
rect 7285 1235 7343 1241
rect 8662 1232 8668 1244
rect 8720 1232 8726 1284
rect 8938 1232 8944 1284
rect 8996 1272 9002 1284
rect 9309 1275 9367 1281
rect 9309 1272 9321 1275
rect 8996 1244 9321 1272
rect 8996 1232 9002 1244
rect 9309 1241 9321 1244
rect 9355 1241 9367 1275
rect 9858 1272 9864 1284
rect 9819 1244 9864 1272
rect 9309 1235 9367 1241
rect 9858 1232 9864 1244
rect 9916 1232 9922 1284
rect 10077 1275 10135 1281
rect 10077 1241 10089 1275
rect 10123 1272 10135 1275
rect 10502 1272 10508 1284
rect 10123 1244 10508 1272
rect 10123 1241 10135 1244
rect 10077 1235 10135 1241
rect 10502 1232 10508 1244
rect 10560 1232 10566 1284
rect 7650 1204 7656 1216
rect 4816 1176 7656 1204
rect 7650 1164 7656 1176
rect 7708 1164 7714 1216
rect 7745 1207 7803 1213
rect 7745 1173 7757 1207
rect 7791 1204 7803 1207
rect 8110 1204 8116 1216
rect 7791 1176 8116 1204
rect 7791 1173 7803 1176
rect 7745 1167 7803 1173
rect 8110 1164 8116 1176
rect 8168 1164 8174 1216
rect 10226 1204 10232 1216
rect 10187 1176 10232 1204
rect 10226 1164 10232 1176
rect 10284 1164 10290 1216
rect 10612 1204 10640 1312
rect 10781 1309 10793 1343
rect 10827 1340 10839 1343
rect 11238 1340 11244 1352
rect 10827 1312 11244 1340
rect 10827 1309 10839 1312
rect 10781 1303 10839 1309
rect 11238 1300 11244 1312
rect 11296 1300 11302 1352
rect 11330 1300 11336 1352
rect 11388 1340 11394 1352
rect 11388 1312 11560 1340
rect 11388 1300 11394 1312
rect 11422 1272 11428 1284
rect 10796 1244 11428 1272
rect 10796 1204 10824 1244
rect 11422 1232 11428 1244
rect 11480 1232 11486 1284
rect 11532 1281 11560 1312
rect 11606 1300 11612 1352
rect 11664 1340 11670 1352
rect 12345 1343 12403 1349
rect 12345 1340 12357 1343
rect 11664 1312 12357 1340
rect 11664 1300 11670 1312
rect 12345 1309 12357 1312
rect 12391 1340 12403 1343
rect 12550 1340 12578 1380
rect 12391 1312 12578 1340
rect 12621 1343 12679 1349
rect 12391 1309 12403 1312
rect 12345 1303 12403 1309
rect 12621 1309 12633 1343
rect 12667 1309 12679 1343
rect 12728 1340 12756 1380
rect 13630 1368 13636 1380
rect 13688 1368 13694 1420
rect 13173 1343 13231 1349
rect 13173 1340 13185 1343
rect 12728 1312 13185 1340
rect 12621 1303 12679 1309
rect 13173 1309 13185 1312
rect 13219 1309 13231 1343
rect 13173 1303 13231 1309
rect 11517 1275 11575 1281
rect 11517 1241 11529 1275
rect 11563 1241 11575 1275
rect 12066 1272 12072 1284
rect 11517 1235 11575 1241
rect 11624 1244 12072 1272
rect 10612 1176 10824 1204
rect 10873 1207 10931 1213
rect 10873 1173 10885 1207
rect 10919 1204 10931 1207
rect 11624 1204 11652 1244
rect 12066 1232 12072 1244
rect 12124 1272 12130 1284
rect 12636 1272 12664 1303
rect 13262 1300 13268 1352
rect 13320 1340 13326 1352
rect 13449 1343 13507 1349
rect 13449 1340 13461 1343
rect 13320 1312 13461 1340
rect 13320 1300 13326 1312
rect 13449 1309 13461 1312
rect 13495 1340 13507 1343
rect 13722 1340 13728 1352
rect 13495 1312 13728 1340
rect 13495 1309 13507 1312
rect 13449 1303 13507 1309
rect 13722 1300 13728 1312
rect 13780 1300 13786 1352
rect 14274 1300 14280 1352
rect 14332 1340 14338 1352
rect 15013 1343 15071 1349
rect 15013 1340 15025 1343
rect 14332 1312 15025 1340
rect 14332 1300 14338 1312
rect 15013 1309 15025 1312
rect 15059 1309 15071 1343
rect 15838 1340 15844 1352
rect 15799 1312 15844 1340
rect 15013 1303 15071 1309
rect 15838 1300 15844 1312
rect 15896 1300 15902 1352
rect 13078 1272 13084 1284
rect 12124 1244 13084 1272
rect 12124 1232 12130 1244
rect 13078 1232 13084 1244
rect 13136 1232 13142 1284
rect 13906 1272 13912 1284
rect 13188 1244 13912 1272
rect 10919 1176 11652 1204
rect 10919 1173 10931 1176
rect 10873 1167 10931 1173
rect 11698 1164 11704 1216
rect 11756 1213 11762 1216
rect 11756 1207 11775 1213
rect 11763 1173 11775 1207
rect 11756 1167 11775 1173
rect 11885 1207 11943 1213
rect 11885 1173 11897 1207
rect 11931 1204 11943 1207
rect 13188 1204 13216 1244
rect 13906 1232 13912 1244
rect 13964 1232 13970 1284
rect 14090 1272 14096 1284
rect 14051 1244 14096 1272
rect 14090 1232 14096 1244
rect 14148 1232 14154 1284
rect 11931 1176 13216 1204
rect 11931 1173 11943 1176
rect 11885 1167 11943 1173
rect 11756 1164 11762 1167
rect 13262 1164 13268 1216
rect 13320 1204 13326 1216
rect 14293 1207 14351 1213
rect 14293 1204 14305 1207
rect 13320 1176 14305 1204
rect 13320 1164 13326 1176
rect 14293 1173 14305 1176
rect 14339 1173 14351 1207
rect 15654 1204 15660 1216
rect 15615 1176 15660 1204
rect 14293 1167 14351 1173
rect 15654 1164 15660 1176
rect 15712 1164 15718 1216
rect 1104 1114 16836 1136
rect 1104 1062 4898 1114
rect 4950 1062 4962 1114
rect 5014 1062 5026 1114
rect 5078 1062 5090 1114
rect 5142 1062 5154 1114
rect 5206 1062 8846 1114
rect 8898 1062 8910 1114
rect 8962 1062 8974 1114
rect 9026 1062 9038 1114
rect 9090 1062 9102 1114
rect 9154 1062 12794 1114
rect 12846 1062 12858 1114
rect 12910 1062 12922 1114
rect 12974 1062 12986 1114
rect 13038 1062 13050 1114
rect 13102 1062 16836 1114
rect 1104 1040 16836 1062
rect 1210 960 1216 1012
rect 1268 1000 1274 1012
rect 10410 1000 10416 1012
rect 1268 972 10416 1000
rect 1268 960 1274 972
rect 10410 960 10416 972
rect 10468 960 10474 1012
rect 10502 960 10508 1012
rect 10560 1000 10566 1012
rect 14458 1000 14464 1012
rect 10560 972 14464 1000
rect 10560 960 10566 972
rect 14458 960 14464 972
rect 14516 960 14522 1012
rect 474 892 480 944
rect 532 932 538 944
rect 8386 932 8392 944
rect 532 904 8392 932
rect 532 892 538 904
rect 8386 892 8392 904
rect 8444 892 8450 944
rect 9858 892 9864 944
rect 9916 932 9922 944
rect 13998 932 14004 944
rect 9916 904 14004 932
rect 9916 892 9922 904
rect 13998 892 14004 904
rect 14056 892 14062 944
rect 4614 824 4620 876
rect 4672 864 4678 876
rect 16666 864 16672 876
rect 4672 836 16672 864
rect 4672 824 4678 836
rect 16666 824 16672 836
rect 16724 824 16730 876
rect 2774 756 2780 808
rect 2832 796 2838 808
rect 8478 796 8484 808
rect 2832 768 8484 796
rect 2832 756 2838 768
rect 8478 756 8484 768
rect 8536 756 8542 808
rect 9582 756 9588 808
rect 9640 796 9646 808
rect 15838 796 15844 808
rect 9640 768 15844 796
rect 9640 756 9646 768
rect 15838 756 15844 768
rect 15896 756 15902 808
rect 2314 688 2320 740
rect 2372 728 2378 740
rect 2372 700 2774 728
rect 2372 688 2378 700
rect 2746 660 2774 700
rect 5258 688 5264 740
rect 5316 728 5322 740
rect 10318 728 10324 740
rect 5316 700 10324 728
rect 5316 688 5322 700
rect 10318 688 10324 700
rect 10376 688 10382 740
rect 9674 660 9680 672
rect 2746 632 9680 660
rect 9674 620 9680 632
rect 9732 620 9738 672
rect 10226 620 10232 672
rect 10284 660 10290 672
rect 16850 660 16856 672
rect 10284 632 16856 660
rect 10284 620 10290 632
rect 16850 620 16856 632
rect 16908 620 16914 672
rect 6638 552 6644 604
rect 6696 592 6702 604
rect 10686 592 10692 604
rect 6696 564 10692 592
rect 6696 552 6702 564
rect 10686 552 10692 564
rect 10744 552 10750 604
rect 3970 484 3976 536
rect 4028 524 4034 536
rect 11698 524 11704 536
rect 4028 496 11704 524
rect 4028 484 4034 496
rect 11698 484 11704 496
rect 11756 524 11762 536
rect 13354 524 13360 536
rect 11756 496 13360 524
rect 11756 484 11762 496
rect 13354 484 13360 496
rect 13412 484 13418 536
rect 4430 416 4436 468
rect 4488 456 4494 468
rect 11330 456 11336 468
rect 4488 428 11336 456
rect 4488 416 4494 428
rect 11330 416 11336 428
rect 11388 416 11394 468
rect 6362 348 6368 400
rect 6420 388 6426 400
rect 9398 388 9404 400
rect 6420 360 9404 388
rect 6420 348 6426 360
rect 9398 348 9404 360
rect 9456 388 9462 400
rect 16022 388 16028 400
rect 9456 360 16028 388
rect 9456 348 9462 360
rect 16022 348 16028 360
rect 16080 348 16086 400
rect 3234 280 3240 332
rect 3292 320 3298 332
rect 13814 320 13820 332
rect 3292 292 13820 320
rect 3292 280 3298 292
rect 13814 280 13820 292
rect 13872 280 13878 332
rect 2222 212 2228 264
rect 2280 252 2286 264
rect 9858 252 9864 264
rect 2280 224 9864 252
rect 2280 212 2286 224
rect 9858 212 9864 224
rect 9916 212 9922 264
rect 3142 144 3148 196
rect 3200 184 3206 196
rect 11974 184 11980 196
rect 3200 156 11980 184
rect 3200 144 3206 156
rect 11974 144 11980 156
rect 12032 144 12038 196
rect 7742 8 7748 60
rect 7800 48 7806 60
rect 15654 48 15660 60
rect 7800 20 15660 48
rect 7800 8 7806 20
rect 15654 8 15660 20
rect 15712 8 15718 60
<< via1 >>
rect 4898 22822 4950 22874
rect 4962 22822 5014 22874
rect 5026 22822 5078 22874
rect 5090 22822 5142 22874
rect 5154 22822 5206 22874
rect 8846 22822 8898 22874
rect 8910 22822 8962 22874
rect 8974 22822 9026 22874
rect 9038 22822 9090 22874
rect 9102 22822 9154 22874
rect 12794 22822 12846 22874
rect 12858 22822 12910 22874
rect 12922 22822 12974 22874
rect 12986 22822 13038 22874
rect 13050 22822 13102 22874
rect 14188 22584 14240 22636
rect 1492 22491 1544 22500
rect 1492 22457 1501 22491
rect 1501 22457 1535 22491
rect 1535 22457 1544 22491
rect 1492 22448 1544 22457
rect 16948 22380 17000 22432
rect 2924 22278 2976 22330
rect 2988 22278 3040 22330
rect 3052 22278 3104 22330
rect 3116 22278 3168 22330
rect 3180 22278 3232 22330
rect 6872 22278 6924 22330
rect 6936 22278 6988 22330
rect 7000 22278 7052 22330
rect 7064 22278 7116 22330
rect 7128 22278 7180 22330
rect 10820 22278 10872 22330
rect 10884 22278 10936 22330
rect 10948 22278 11000 22330
rect 11012 22278 11064 22330
rect 11076 22278 11128 22330
rect 14768 22278 14820 22330
rect 14832 22278 14884 22330
rect 14896 22278 14948 22330
rect 14960 22278 15012 22330
rect 15024 22278 15076 22330
rect 1584 22219 1636 22228
rect 1584 22185 1593 22219
rect 1593 22185 1627 22219
rect 1627 22185 1636 22219
rect 1584 22176 1636 22185
rect 2780 22151 2832 22160
rect 2780 22117 2789 22151
rect 2789 22117 2823 22151
rect 2823 22117 2832 22151
rect 2780 22108 2832 22117
rect 8024 22040 8076 22092
rect 3884 21972 3936 22024
rect 8576 21904 8628 21956
rect 6736 21836 6788 21888
rect 4898 21734 4950 21786
rect 4962 21734 5014 21786
rect 5026 21734 5078 21786
rect 5090 21734 5142 21786
rect 5154 21734 5206 21786
rect 8846 21734 8898 21786
rect 8910 21734 8962 21786
rect 8974 21734 9026 21786
rect 9038 21734 9090 21786
rect 9102 21734 9154 21786
rect 12794 21734 12846 21786
rect 12858 21734 12910 21786
rect 12922 21734 12974 21786
rect 12986 21734 13038 21786
rect 13050 21734 13102 21786
rect 388 21632 440 21684
rect 4068 21428 4120 21480
rect 9312 21360 9364 21412
rect 1400 21292 1452 21344
rect 3424 21292 3476 21344
rect 3608 21335 3660 21344
rect 3608 21301 3617 21335
rect 3617 21301 3651 21335
rect 3651 21301 3660 21335
rect 3608 21292 3660 21301
rect 2924 21190 2976 21242
rect 2988 21190 3040 21242
rect 3052 21190 3104 21242
rect 3116 21190 3168 21242
rect 3180 21190 3232 21242
rect 6872 21190 6924 21242
rect 6936 21190 6988 21242
rect 7000 21190 7052 21242
rect 7064 21190 7116 21242
rect 7128 21190 7180 21242
rect 10820 21190 10872 21242
rect 10884 21190 10936 21242
rect 10948 21190 11000 21242
rect 11012 21190 11064 21242
rect 11076 21190 11128 21242
rect 14768 21190 14820 21242
rect 14832 21190 14884 21242
rect 14896 21190 14948 21242
rect 14960 21190 15012 21242
rect 15024 21190 15076 21242
rect 2412 21131 2464 21140
rect 2412 21097 2421 21131
rect 2421 21097 2455 21131
rect 2455 21097 2464 21131
rect 2412 21088 2464 21097
rect 1492 20927 1544 20936
rect 1492 20893 1501 20927
rect 1501 20893 1535 20927
rect 1535 20893 1544 20927
rect 1492 20884 1544 20893
rect 2228 20927 2280 20936
rect 2228 20893 2237 20927
rect 2237 20893 2271 20927
rect 2271 20893 2280 20927
rect 2228 20884 2280 20893
rect 2780 20884 2832 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 10416 20884 10468 20936
rect 2688 20816 2740 20868
rect 3608 20816 3660 20868
rect 1584 20748 1636 20800
rect 3700 20748 3752 20800
rect 3792 20791 3844 20800
rect 3792 20757 3801 20791
rect 3801 20757 3835 20791
rect 3835 20757 3844 20791
rect 3792 20748 3844 20757
rect 4160 20748 4212 20800
rect 4898 20646 4950 20698
rect 4962 20646 5014 20698
rect 5026 20646 5078 20698
rect 5090 20646 5142 20698
rect 5154 20646 5206 20698
rect 8846 20646 8898 20698
rect 8910 20646 8962 20698
rect 8974 20646 9026 20698
rect 9038 20646 9090 20698
rect 9102 20646 9154 20698
rect 12794 20646 12846 20698
rect 12858 20646 12910 20698
rect 12922 20646 12974 20698
rect 12986 20646 13038 20698
rect 13050 20646 13102 20698
rect 2780 20544 2832 20596
rect 4620 20544 4672 20596
rect 1032 20408 1084 20460
rect 3148 20408 3200 20460
rect 4160 20408 4212 20460
rect 4252 20451 4304 20460
rect 4252 20417 4261 20451
rect 4261 20417 4295 20451
rect 4295 20417 4304 20451
rect 15292 20476 15344 20528
rect 4252 20408 4304 20417
rect 3332 20340 3384 20392
rect 9680 20408 9732 20460
rect 17316 20408 17368 20460
rect 2412 20272 2464 20324
rect 3516 20272 3568 20324
rect 4160 20272 4212 20324
rect 16028 20272 16080 20324
rect 1768 20204 1820 20256
rect 1860 20204 1912 20256
rect 2320 20204 2372 20256
rect 4804 20204 4856 20256
rect 5724 20204 5776 20256
rect 5816 20204 5868 20256
rect 17408 20204 17460 20256
rect 2924 20102 2976 20154
rect 2988 20102 3040 20154
rect 3052 20102 3104 20154
rect 3116 20102 3168 20154
rect 3180 20102 3232 20154
rect 6872 20102 6924 20154
rect 6936 20102 6988 20154
rect 7000 20102 7052 20154
rect 7064 20102 7116 20154
rect 7128 20102 7180 20154
rect 10820 20102 10872 20154
rect 10884 20102 10936 20154
rect 10948 20102 11000 20154
rect 11012 20102 11064 20154
rect 11076 20102 11128 20154
rect 14768 20102 14820 20154
rect 14832 20102 14884 20154
rect 14896 20102 14948 20154
rect 14960 20102 15012 20154
rect 15024 20102 15076 20154
rect 3976 20000 4028 20052
rect 4804 20000 4856 20052
rect 17224 20000 17276 20052
rect 3516 19932 3568 19984
rect 3792 19975 3844 19984
rect 3792 19941 3801 19975
rect 3801 19941 3835 19975
rect 3835 19941 3844 19975
rect 3792 19932 3844 19941
rect 5356 19975 5408 19984
rect 5356 19941 5365 19975
rect 5365 19941 5399 19975
rect 5399 19941 5408 19975
rect 5356 19932 5408 19941
rect 3608 19864 3660 19916
rect 2872 19728 2924 19780
rect 3332 19796 3384 19848
rect 4160 19864 4212 19916
rect 4344 19796 4396 19848
rect 4528 19839 4580 19848
rect 4528 19805 4537 19839
rect 4537 19805 4571 19839
rect 4571 19805 4580 19839
rect 4528 19796 4580 19805
rect 6460 19864 6512 19916
rect 5816 19839 5868 19848
rect 5816 19805 5825 19839
rect 5825 19805 5859 19839
rect 5859 19805 5868 19839
rect 5816 19796 5868 19805
rect 3516 19728 3568 19780
rect 3608 19660 3660 19712
rect 3976 19660 4028 19712
rect 4344 19660 4396 19712
rect 5632 19728 5684 19780
rect 5816 19660 5868 19712
rect 6000 19660 6052 19712
rect 12532 19796 12584 19848
rect 14004 19660 14056 19712
rect 4898 19558 4950 19610
rect 4962 19558 5014 19610
rect 5026 19558 5078 19610
rect 5090 19558 5142 19610
rect 5154 19558 5206 19610
rect 8846 19558 8898 19610
rect 8910 19558 8962 19610
rect 8974 19558 9026 19610
rect 9038 19558 9090 19610
rect 9102 19558 9154 19610
rect 12794 19558 12846 19610
rect 12858 19558 12910 19610
rect 12922 19558 12974 19610
rect 12986 19558 13038 19610
rect 13050 19558 13102 19610
rect 1492 19456 1544 19508
rect 3148 19456 3200 19508
rect 1492 19320 1544 19372
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 2596 19388 2648 19440
rect 2688 19388 2740 19440
rect 4160 19456 4212 19508
rect 4528 19456 4580 19508
rect 3516 19431 3568 19440
rect 3516 19397 3525 19431
rect 3525 19397 3559 19431
rect 3559 19397 3568 19431
rect 3516 19388 3568 19397
rect 2320 19320 2372 19372
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 5264 19388 5316 19440
rect 5540 19456 5592 19508
rect 6092 19388 6144 19440
rect 15476 19388 15528 19440
rect 2044 19295 2096 19304
rect 2044 19261 2053 19295
rect 2053 19261 2087 19295
rect 2087 19261 2096 19295
rect 2044 19252 2096 19261
rect 2596 19252 2648 19304
rect 5264 19252 5316 19304
rect 3148 19184 3200 19236
rect 4804 19116 4856 19168
rect 5908 19184 5960 19236
rect 6644 19320 6696 19372
rect 10692 19320 10744 19372
rect 7472 19184 7524 19236
rect 5172 19116 5224 19168
rect 5816 19116 5868 19168
rect 17592 19184 17644 19236
rect 2924 19014 2976 19066
rect 2988 19014 3040 19066
rect 3052 19014 3104 19066
rect 3116 19014 3168 19066
rect 3180 19014 3232 19066
rect 6872 19014 6924 19066
rect 6936 19014 6988 19066
rect 7000 19014 7052 19066
rect 7064 19014 7116 19066
rect 7128 19014 7180 19066
rect 10820 19014 10872 19066
rect 10884 19014 10936 19066
rect 10948 19014 11000 19066
rect 11012 19014 11064 19066
rect 11076 19014 11128 19066
rect 14768 19014 14820 19066
rect 14832 19014 14884 19066
rect 14896 19014 14948 19066
rect 14960 19014 15012 19066
rect 15024 19014 15076 19066
rect 2780 18844 2832 18896
rect 4712 18912 4764 18964
rect 3056 18819 3108 18828
rect 3056 18785 3065 18819
rect 3065 18785 3099 18819
rect 3099 18785 3108 18819
rect 3056 18776 3108 18785
rect 3884 18844 3936 18896
rect 3976 18844 4028 18896
rect 8300 18912 8352 18964
rect 2320 18708 2372 18760
rect 5724 18751 5776 18760
rect 5724 18717 5733 18751
rect 5733 18717 5767 18751
rect 5767 18717 5776 18751
rect 5724 18708 5776 18717
rect 6092 18776 6144 18828
rect 13912 18912 13964 18964
rect 8484 18844 8536 18896
rect 13452 18844 13504 18896
rect 6184 18751 6236 18760
rect 6184 18717 6193 18751
rect 6193 18717 6227 18751
rect 6227 18717 6236 18751
rect 6184 18708 6236 18717
rect 8760 18776 8812 18828
rect 13820 18776 13872 18828
rect 6552 18751 6604 18760
rect 6552 18717 6561 18751
rect 6561 18717 6595 18751
rect 6595 18717 6604 18751
rect 7104 18751 7156 18760
rect 6552 18708 6604 18717
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 17040 18708 17092 18760
rect 2780 18640 2832 18692
rect 2596 18572 2648 18624
rect 3792 18640 3844 18692
rect 4068 18640 4120 18692
rect 16856 18640 16908 18692
rect 3884 18572 3936 18624
rect 4528 18572 4580 18624
rect 5816 18572 5868 18624
rect 8300 18572 8352 18624
rect 10784 18572 10836 18624
rect 4898 18470 4950 18522
rect 4962 18470 5014 18522
rect 5026 18470 5078 18522
rect 5090 18470 5142 18522
rect 5154 18470 5206 18522
rect 8846 18470 8898 18522
rect 8910 18470 8962 18522
rect 8974 18470 9026 18522
rect 9038 18470 9090 18522
rect 9102 18470 9154 18522
rect 12794 18470 12846 18522
rect 12858 18470 12910 18522
rect 12922 18470 12974 18522
rect 12986 18470 13038 18522
rect 13050 18470 13102 18522
rect 1952 18368 2004 18420
rect 3240 18368 3292 18420
rect 1308 18300 1360 18352
rect 6276 18368 6328 18420
rect 7472 18411 7524 18420
rect 7472 18377 7481 18411
rect 7481 18377 7515 18411
rect 7515 18377 7524 18411
rect 7472 18368 7524 18377
rect 8576 18368 8628 18420
rect 9036 18368 9088 18420
rect 9312 18368 9364 18420
rect 9496 18411 9548 18420
rect 9496 18377 9505 18411
rect 9505 18377 9539 18411
rect 9539 18377 9548 18411
rect 9496 18368 9548 18377
rect 1768 18232 1820 18284
rect 2872 18232 2924 18284
rect 3700 18232 3752 18284
rect 6460 18300 6512 18352
rect 9956 18300 10008 18352
rect 7196 18232 7248 18284
rect 8024 18275 8076 18284
rect 8024 18241 8033 18275
rect 8033 18241 8067 18275
rect 8067 18241 8076 18275
rect 8024 18232 8076 18241
rect 8300 18232 8352 18284
rect 3792 18207 3844 18216
rect 3792 18173 3801 18207
rect 3801 18173 3835 18207
rect 3835 18173 3844 18207
rect 3792 18164 3844 18173
rect 7472 18164 7524 18216
rect 16212 18232 16264 18284
rect 11796 18164 11848 18216
rect 3424 18028 3476 18080
rect 4068 18028 4120 18080
rect 12440 18096 12492 18148
rect 5172 18071 5224 18080
rect 5172 18037 5181 18071
rect 5181 18037 5215 18071
rect 5215 18037 5224 18071
rect 5172 18028 5224 18037
rect 6276 18028 6328 18080
rect 8116 18028 8168 18080
rect 8760 18028 8812 18080
rect 17132 18028 17184 18080
rect 2924 17926 2976 17978
rect 2988 17926 3040 17978
rect 3052 17926 3104 17978
rect 3116 17926 3168 17978
rect 3180 17926 3232 17978
rect 6872 17926 6924 17978
rect 6936 17926 6988 17978
rect 7000 17926 7052 17978
rect 7064 17926 7116 17978
rect 7128 17926 7180 17978
rect 10820 17926 10872 17978
rect 10884 17926 10936 17978
rect 10948 17926 11000 17978
rect 11012 17926 11064 17978
rect 11076 17926 11128 17978
rect 14768 17926 14820 17978
rect 14832 17926 14884 17978
rect 14896 17926 14948 17978
rect 14960 17926 15012 17978
rect 15024 17926 15076 17978
rect 296 17824 348 17876
rect 5724 17824 5776 17876
rect 6276 17824 6328 17876
rect 9312 17824 9364 17876
rect 8024 17756 8076 17808
rect 8392 17756 8444 17808
rect 10692 17824 10744 17876
rect 15384 17824 15436 17876
rect 9588 17756 9640 17808
rect 1952 17620 2004 17672
rect 1124 17552 1176 17604
rect 2596 17552 2648 17604
rect 4160 17620 4212 17672
rect 6092 17688 6144 17740
rect 7472 17688 7524 17740
rect 8576 17688 8628 17740
rect 9220 17688 9272 17740
rect 3700 17484 3752 17536
rect 4712 17552 4764 17604
rect 6552 17552 6604 17604
rect 5816 17484 5868 17536
rect 7380 17620 7432 17672
rect 7748 17620 7800 17672
rect 8116 17620 8168 17672
rect 9128 17663 9180 17672
rect 7104 17595 7156 17604
rect 7104 17561 7113 17595
rect 7113 17561 7147 17595
rect 7147 17561 7156 17595
rect 7104 17552 7156 17561
rect 7840 17552 7892 17604
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 9588 17663 9640 17672
rect 9588 17629 9597 17663
rect 9597 17629 9631 17663
rect 9631 17629 9640 17663
rect 9588 17620 9640 17629
rect 10140 17620 10192 17672
rect 8484 17552 8536 17604
rect 8576 17552 8628 17604
rect 9036 17552 9088 17604
rect 9312 17552 9364 17604
rect 9496 17552 9548 17604
rect 15660 17552 15712 17604
rect 8852 17484 8904 17536
rect 10048 17484 10100 17536
rect 10232 17484 10284 17536
rect 14464 17484 14516 17536
rect 4898 17382 4950 17434
rect 4962 17382 5014 17434
rect 5026 17382 5078 17434
rect 5090 17382 5142 17434
rect 5154 17382 5206 17434
rect 8846 17382 8898 17434
rect 8910 17382 8962 17434
rect 8974 17382 9026 17434
rect 9038 17382 9090 17434
rect 9102 17382 9154 17434
rect 12794 17382 12846 17434
rect 12858 17382 12910 17434
rect 12922 17382 12974 17434
rect 12986 17382 13038 17434
rect 13050 17382 13102 17434
rect 6460 17280 6512 17332
rect 2136 17212 2188 17264
rect 1952 17187 2004 17196
rect 1952 17153 1961 17187
rect 1961 17153 1995 17187
rect 1995 17153 2004 17187
rect 1952 17144 2004 17153
rect 2964 17144 3016 17196
rect 3792 17187 3844 17196
rect 3792 17153 3801 17187
rect 3801 17153 3835 17187
rect 3835 17153 3844 17187
rect 3792 17144 3844 17153
rect 6000 17144 6052 17196
rect 6276 17144 6328 17196
rect 10232 17280 10284 17332
rect 10692 17280 10744 17332
rect 13636 17280 13688 17332
rect 7656 17212 7708 17264
rect 15752 17212 15804 17264
rect 7840 17187 7892 17196
rect 6460 17076 6512 17128
rect 7380 17119 7432 17128
rect 7380 17085 7389 17119
rect 7389 17085 7423 17119
rect 7423 17085 7432 17119
rect 7380 17076 7432 17085
rect 5724 17008 5776 17060
rect 7564 17008 7616 17060
rect 7840 17153 7849 17187
rect 7849 17153 7883 17187
rect 7883 17153 7892 17187
rect 7840 17144 7892 17153
rect 7932 17144 7984 17196
rect 9036 17187 9088 17196
rect 9036 17153 9045 17187
rect 9045 17153 9079 17187
rect 9079 17153 9088 17187
rect 9680 17187 9732 17196
rect 9036 17144 9088 17153
rect 7748 17076 7800 17128
rect 8576 17076 8628 17128
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 8024 17008 8076 17060
rect 9404 17008 9456 17060
rect 10324 17076 10376 17128
rect 15108 17076 15160 17128
rect 16764 17008 16816 17060
rect 4436 16940 4488 16992
rect 6000 16940 6052 16992
rect 6644 16940 6696 16992
rect 9680 16940 9732 16992
rect 10508 16940 10560 16992
rect 10600 16940 10652 16992
rect 14280 16940 14332 16992
rect 2924 16838 2976 16890
rect 2988 16838 3040 16890
rect 3052 16838 3104 16890
rect 3116 16838 3168 16890
rect 3180 16838 3232 16890
rect 6872 16838 6924 16890
rect 6936 16838 6988 16890
rect 7000 16838 7052 16890
rect 7064 16838 7116 16890
rect 7128 16838 7180 16890
rect 10820 16838 10872 16890
rect 10884 16838 10936 16890
rect 10948 16838 11000 16890
rect 11012 16838 11064 16890
rect 11076 16838 11128 16890
rect 14768 16838 14820 16890
rect 14832 16838 14884 16890
rect 14896 16838 14948 16890
rect 14960 16838 15012 16890
rect 15024 16838 15076 16890
rect 848 16736 900 16788
rect 6184 16736 6236 16788
rect 7748 16736 7800 16788
rect 8024 16736 8076 16788
rect 8300 16736 8352 16788
rect 9496 16736 9548 16788
rect 9772 16736 9824 16788
rect 10324 16736 10376 16788
rect 5448 16668 5500 16720
rect 2596 16532 2648 16584
rect 4528 16575 4580 16584
rect 4528 16541 4537 16575
rect 4537 16541 4571 16575
rect 4571 16541 4580 16575
rect 6368 16600 6420 16652
rect 8944 16668 8996 16720
rect 10784 16736 10836 16788
rect 16580 16736 16632 16788
rect 4528 16532 4580 16541
rect 8300 16532 8352 16584
rect 8576 16532 8628 16584
rect 10600 16600 10652 16652
rect 8944 16532 8996 16584
rect 9128 16532 9180 16584
rect 11704 16575 11756 16584
rect 11704 16541 11713 16575
rect 11713 16541 11747 16575
rect 11747 16541 11756 16575
rect 11704 16532 11756 16541
rect 1768 16464 1820 16516
rect 756 16396 808 16448
rect 1492 16396 1544 16448
rect 3332 16396 3384 16448
rect 4068 16464 4120 16516
rect 7104 16464 7156 16516
rect 4620 16439 4672 16448
rect 4620 16405 4629 16439
rect 4629 16405 4663 16439
rect 4663 16405 4672 16439
rect 4620 16396 4672 16405
rect 4804 16439 4856 16448
rect 4804 16405 4813 16439
rect 4813 16405 4847 16439
rect 4847 16405 4856 16439
rect 4804 16396 4856 16405
rect 5540 16396 5592 16448
rect 6368 16396 6420 16448
rect 6828 16396 6880 16448
rect 7288 16396 7340 16448
rect 7380 16396 7432 16448
rect 8208 16396 8260 16448
rect 8484 16396 8536 16448
rect 8668 16464 8720 16516
rect 9220 16464 9272 16516
rect 9680 16396 9732 16448
rect 9864 16396 9916 16448
rect 10876 16396 10928 16448
rect 14556 16464 14608 16516
rect 4898 16294 4950 16346
rect 4962 16294 5014 16346
rect 5026 16294 5078 16346
rect 5090 16294 5142 16346
rect 5154 16294 5206 16346
rect 8846 16294 8898 16346
rect 8910 16294 8962 16346
rect 8974 16294 9026 16346
rect 9038 16294 9090 16346
rect 9102 16294 9154 16346
rect 12794 16294 12846 16346
rect 12858 16294 12910 16346
rect 12922 16294 12974 16346
rect 12986 16294 13038 16346
rect 13050 16294 13102 16346
rect 2228 16192 2280 16244
rect 2412 16192 2464 16244
rect 2688 16192 2740 16244
rect 1216 16056 1268 16108
rect 2504 16124 2556 16176
rect 2872 16167 2924 16176
rect 2872 16133 2906 16167
rect 2906 16133 2924 16167
rect 2872 16124 2924 16133
rect 3976 16124 4028 16176
rect 4528 16124 4580 16176
rect 8024 16192 8076 16244
rect 5908 16124 5960 16176
rect 8300 16192 8352 16244
rect 8760 16192 8812 16244
rect 8484 16124 8536 16176
rect 9772 16192 9824 16244
rect 10600 16192 10652 16244
rect 9404 16124 9456 16176
rect 2228 16056 2280 16108
rect 6184 16056 6236 16108
rect 6644 16099 6696 16108
rect 6644 16065 6653 16099
rect 6653 16065 6687 16099
rect 6687 16065 6696 16099
rect 6644 16056 6696 16065
rect 6736 16056 6788 16108
rect 7196 16099 7248 16108
rect 7196 16065 7205 16099
rect 7205 16065 7239 16099
rect 7239 16065 7248 16099
rect 7196 16056 7248 16065
rect 7932 16099 7984 16108
rect 7932 16065 7941 16099
rect 7941 16065 7975 16099
rect 7975 16065 7984 16099
rect 7932 16056 7984 16065
rect 8116 16099 8168 16108
rect 8116 16065 8125 16099
rect 8125 16065 8159 16099
rect 8159 16065 8168 16099
rect 8116 16056 8168 16065
rect 8300 16099 8352 16108
rect 8300 16065 8309 16099
rect 8309 16065 8343 16099
rect 8343 16065 8352 16099
rect 8300 16056 8352 16065
rect 9588 16056 9640 16108
rect 9864 16099 9916 16108
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 1860 16031 1912 16040
rect 1860 15997 1869 16031
rect 1869 15997 1903 16031
rect 1903 15997 1912 16031
rect 1860 15988 1912 15997
rect 2596 16031 2648 16040
rect 2596 15997 2605 16031
rect 2605 15997 2639 16031
rect 2639 15997 2648 16031
rect 2596 15988 2648 15997
rect 3700 15852 3752 15904
rect 5908 15920 5960 15972
rect 9312 15988 9364 16040
rect 9864 16065 9873 16099
rect 9873 16065 9907 16099
rect 9907 16065 9916 16099
rect 9864 16056 9916 16065
rect 10232 16124 10284 16176
rect 12164 16192 12216 16244
rect 14096 16124 14148 16176
rect 10600 16099 10652 16108
rect 10600 16065 10609 16099
rect 10609 16065 10643 16099
rect 10643 16065 10652 16099
rect 10600 16056 10652 16065
rect 10876 16099 10928 16108
rect 10876 16065 10885 16099
rect 10885 16065 10919 16099
rect 10919 16065 10928 16099
rect 10876 16056 10928 16065
rect 11612 16056 11664 16108
rect 11244 15988 11296 16040
rect 11888 16056 11940 16108
rect 15292 16056 15344 16108
rect 16488 16056 16540 16108
rect 7104 15920 7156 15972
rect 8668 15920 8720 15972
rect 8852 15920 8904 15972
rect 5724 15852 5776 15904
rect 6368 15852 6420 15904
rect 6644 15852 6696 15904
rect 6828 15852 6880 15904
rect 6920 15852 6972 15904
rect 8300 15852 8352 15904
rect 8760 15852 8812 15904
rect 9588 15852 9640 15904
rect 9864 15920 9916 15972
rect 12624 15920 12676 15972
rect 15292 15920 15344 15972
rect 9956 15852 10008 15904
rect 10692 15852 10744 15904
rect 10784 15852 10836 15904
rect 11336 15852 11388 15904
rect 11520 15895 11572 15904
rect 11520 15861 11529 15895
rect 11529 15861 11563 15895
rect 11563 15861 11572 15895
rect 11520 15852 11572 15861
rect 11704 15852 11756 15904
rect 2924 15750 2976 15802
rect 2988 15750 3040 15802
rect 3052 15750 3104 15802
rect 3116 15750 3168 15802
rect 3180 15750 3232 15802
rect 6872 15750 6924 15802
rect 6936 15750 6988 15802
rect 7000 15750 7052 15802
rect 7064 15750 7116 15802
rect 7128 15750 7180 15802
rect 10820 15750 10872 15802
rect 10884 15750 10936 15802
rect 10948 15750 11000 15802
rect 11012 15750 11064 15802
rect 11076 15750 11128 15802
rect 14768 15750 14820 15802
rect 14832 15750 14884 15802
rect 14896 15750 14948 15802
rect 14960 15750 15012 15802
rect 15024 15750 15076 15802
rect 2136 15648 2188 15700
rect 3976 15691 4028 15700
rect 3976 15657 3985 15691
rect 3985 15657 4019 15691
rect 4019 15657 4028 15691
rect 3976 15648 4028 15657
rect 5632 15648 5684 15700
rect 6552 15691 6604 15700
rect 6552 15657 6561 15691
rect 6561 15657 6595 15691
rect 6595 15657 6604 15691
rect 6552 15648 6604 15657
rect 1400 15580 1452 15632
rect 2596 15580 2648 15632
rect 3792 15580 3844 15632
rect 4160 15580 4212 15632
rect 2504 15512 2556 15564
rect 12164 15648 12216 15700
rect 13084 15691 13136 15700
rect 13084 15657 13093 15691
rect 13093 15657 13127 15691
rect 13127 15657 13136 15691
rect 13084 15648 13136 15657
rect 14556 15691 14608 15700
rect 14556 15657 14565 15691
rect 14565 15657 14599 15691
rect 14599 15657 14608 15691
rect 14556 15648 14608 15657
rect 7748 15580 7800 15632
rect 8300 15512 8352 15564
rect 9496 15512 9548 15564
rect 3792 15444 3844 15496
rect 2320 15376 2372 15428
rect 4344 15376 4396 15428
rect 1400 15308 1452 15360
rect 3976 15308 4028 15360
rect 5540 15444 5592 15496
rect 8484 15444 8536 15496
rect 9036 15444 9088 15496
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 10048 15487 10100 15496
rect 9404 15444 9456 15453
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 10968 15580 11020 15632
rect 11336 15580 11388 15632
rect 12532 15580 12584 15632
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 12256 15512 12308 15564
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10784 15487 10836 15496
rect 10324 15444 10376 15453
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 10784 15444 10836 15453
rect 5080 15308 5132 15360
rect 6092 15308 6144 15360
rect 8668 15308 8720 15360
rect 8944 15351 8996 15360
rect 8944 15317 8953 15351
rect 8953 15317 8987 15351
rect 8987 15317 8996 15351
rect 8944 15308 8996 15317
rect 9220 15308 9272 15360
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 10048 15308 10100 15360
rect 10600 15376 10652 15428
rect 11428 15444 11480 15496
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 12900 15512 12952 15564
rect 12992 15487 13044 15496
rect 12992 15453 13001 15487
rect 13001 15453 13035 15487
rect 13035 15453 13044 15487
rect 12992 15444 13044 15453
rect 11520 15308 11572 15360
rect 11704 15308 11756 15360
rect 11980 15308 12032 15360
rect 13360 15376 13412 15428
rect 15844 15444 15896 15496
rect 16672 15308 16724 15360
rect 4898 15206 4950 15258
rect 4962 15206 5014 15258
rect 5026 15206 5078 15258
rect 5090 15206 5142 15258
rect 5154 15206 5206 15258
rect 8846 15206 8898 15258
rect 8910 15206 8962 15258
rect 8974 15206 9026 15258
rect 9038 15206 9090 15258
rect 9102 15206 9154 15258
rect 12794 15206 12846 15258
rect 12858 15206 12910 15258
rect 12922 15206 12974 15258
rect 12986 15206 13038 15258
rect 13050 15206 13102 15258
rect 1860 15104 1912 15156
rect 2228 15104 2280 15156
rect 4528 15104 4580 15156
rect 5356 15104 5408 15156
rect 1584 15011 1636 15020
rect 1584 14977 1602 15011
rect 1602 14977 1636 15011
rect 2688 15036 2740 15088
rect 2964 15036 3016 15088
rect 4620 15036 4672 15088
rect 5908 15036 5960 15088
rect 6276 15036 6328 15088
rect 8300 15104 8352 15156
rect 9036 15104 9088 15156
rect 9312 15104 9364 15156
rect 11336 15104 11388 15156
rect 11704 15147 11756 15156
rect 11704 15113 11713 15147
rect 11713 15113 11747 15147
rect 11747 15113 11756 15147
rect 11704 15104 11756 15113
rect 12256 15104 12308 15156
rect 13544 15104 13596 15156
rect 13728 15104 13780 15156
rect 15660 15147 15712 15156
rect 15660 15113 15669 15147
rect 15669 15113 15703 15147
rect 15703 15113 15712 15147
rect 15660 15104 15712 15113
rect 8116 15036 8168 15088
rect 1860 15011 1912 15020
rect 1584 14968 1636 14977
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 2320 14968 2372 15020
rect 2872 15011 2924 15020
rect 1768 14900 1820 14952
rect 2872 14977 2906 15011
rect 2906 14977 2924 15011
rect 2872 14968 2924 14977
rect 6552 14968 6604 15020
rect 6644 15011 6696 15020
rect 6644 14977 6653 15011
rect 6653 14977 6687 15011
rect 6687 14977 6696 15011
rect 7196 15011 7248 15020
rect 6644 14968 6696 14977
rect 7196 14977 7205 15011
rect 7205 14977 7239 15011
rect 7239 14977 7248 15011
rect 7196 14968 7248 14977
rect 8300 14968 8352 15020
rect 9312 14968 9364 15020
rect 9680 14968 9732 15020
rect 2596 14943 2648 14952
rect 2596 14909 2605 14943
rect 2605 14909 2639 14943
rect 2639 14909 2648 14943
rect 2596 14900 2648 14909
rect 4160 14900 4212 14952
rect 6184 14900 6236 14952
rect 7472 14900 7524 14952
rect 9956 14900 10008 14952
rect 10324 14968 10376 15020
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 11428 15036 11480 15088
rect 15936 15036 15988 15088
rect 11704 14900 11756 14952
rect 12440 15011 12492 15020
rect 12440 14977 12441 15011
rect 12441 14977 12475 15011
rect 12475 14977 12492 15011
rect 12440 14968 12492 14977
rect 12900 14968 12952 15020
rect 13728 15011 13780 15020
rect 13728 14977 13737 15011
rect 13737 14977 13771 15011
rect 13771 14977 13780 15011
rect 13728 14968 13780 14977
rect 13820 14968 13872 15020
rect 15568 15011 15620 15020
rect 15568 14977 15577 15011
rect 15577 14977 15611 15011
rect 15611 14977 15620 15011
rect 15568 14968 15620 14977
rect 14188 14900 14240 14952
rect 1584 14832 1636 14884
rect 5632 14832 5684 14884
rect 10600 14832 10652 14884
rect 1768 14764 1820 14816
rect 4160 14764 4212 14816
rect 5908 14764 5960 14816
rect 8852 14764 8904 14816
rect 8944 14764 8996 14816
rect 9680 14764 9732 14816
rect 15660 14832 15712 14884
rect 11612 14764 11664 14816
rect 12440 14764 12492 14816
rect 13268 14807 13320 14816
rect 13268 14773 13277 14807
rect 13277 14773 13311 14807
rect 13311 14773 13320 14807
rect 13268 14764 13320 14773
rect 2924 14662 2976 14714
rect 2988 14662 3040 14714
rect 3052 14662 3104 14714
rect 3116 14662 3168 14714
rect 3180 14662 3232 14714
rect 6872 14662 6924 14714
rect 6936 14662 6988 14714
rect 7000 14662 7052 14714
rect 7064 14662 7116 14714
rect 7128 14662 7180 14714
rect 10820 14662 10872 14714
rect 10884 14662 10936 14714
rect 10948 14662 11000 14714
rect 11012 14662 11064 14714
rect 11076 14662 11128 14714
rect 14768 14662 14820 14714
rect 14832 14662 14884 14714
rect 14896 14662 14948 14714
rect 14960 14662 15012 14714
rect 15024 14662 15076 14714
rect 1860 14560 1912 14612
rect 1584 14424 1636 14476
rect 7012 14560 7064 14612
rect 7104 14560 7156 14612
rect 7288 14560 7340 14612
rect 5632 14535 5684 14544
rect 5632 14501 5641 14535
rect 5641 14501 5675 14535
rect 5675 14501 5684 14535
rect 5632 14492 5684 14501
rect 5908 14356 5960 14408
rect 7380 14356 7432 14408
rect 7748 14560 7800 14612
rect 8852 14560 8904 14612
rect 11520 14560 11572 14612
rect 1400 14288 1452 14340
rect 1584 14288 1636 14340
rect 6460 14288 6512 14340
rect 6552 14288 6604 14340
rect 8300 14424 8352 14476
rect 8576 14424 8628 14476
rect 8760 14492 8812 14544
rect 9036 14492 9088 14544
rect 9128 14492 9180 14544
rect 10416 14492 10468 14544
rect 10600 14492 10652 14544
rect 12072 14560 12124 14612
rect 12900 14560 12952 14612
rect 14280 14560 14332 14612
rect 8484 14356 8536 14408
rect 9036 14356 9088 14408
rect 9864 14424 9916 14476
rect 10876 14467 10928 14476
rect 10876 14433 10885 14467
rect 10885 14433 10919 14467
rect 10919 14433 10928 14467
rect 10876 14424 10928 14433
rect 11428 14356 11480 14408
rect 1216 14220 1268 14272
rect 1860 14220 1912 14272
rect 2412 14220 2464 14272
rect 8576 14288 8628 14340
rect 8668 14288 8720 14340
rect 9220 14288 9272 14340
rect 9772 14288 9824 14340
rect 11244 14288 11296 14340
rect 11520 14288 11572 14340
rect 12532 14424 12584 14476
rect 12716 14424 12768 14476
rect 13544 14424 13596 14476
rect 12164 14356 12216 14408
rect 13176 14356 13228 14408
rect 13452 14399 13504 14408
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13452 14356 13504 14365
rect 13636 14356 13688 14408
rect 14004 14356 14056 14408
rect 14924 14399 14976 14408
rect 14924 14365 14933 14399
rect 14933 14365 14967 14399
rect 14967 14365 14976 14399
rect 14924 14356 14976 14365
rect 14648 14288 14700 14340
rect 7196 14220 7248 14272
rect 9404 14220 9456 14272
rect 9496 14220 9548 14272
rect 10692 14220 10744 14272
rect 11336 14220 11388 14272
rect 11612 14220 11664 14272
rect 11704 14220 11756 14272
rect 13636 14220 13688 14272
rect 13820 14220 13872 14272
rect 15016 14220 15068 14272
rect 4898 14118 4950 14170
rect 4962 14118 5014 14170
rect 5026 14118 5078 14170
rect 5090 14118 5142 14170
rect 5154 14118 5206 14170
rect 8846 14118 8898 14170
rect 8910 14118 8962 14170
rect 8974 14118 9026 14170
rect 9038 14118 9090 14170
rect 9102 14118 9154 14170
rect 12794 14118 12846 14170
rect 12858 14118 12910 14170
rect 12922 14118 12974 14170
rect 12986 14118 13038 14170
rect 13050 14118 13102 14170
rect 1216 14016 1268 14068
rect 1124 13948 1176 14000
rect 1400 13948 1452 14000
rect 1768 13991 1820 14000
rect 1768 13957 1777 13991
rect 1777 13957 1811 13991
rect 1811 13957 1820 13991
rect 1768 13948 1820 13957
rect 2228 13948 2280 14000
rect 756 13880 808 13932
rect 1768 13812 1820 13864
rect 2412 13880 2464 13932
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 3976 13880 4028 13932
rect 6644 14016 6696 14068
rect 7564 14016 7616 14068
rect 8944 14016 8996 14068
rect 7472 13948 7524 14000
rect 7748 13948 7800 14000
rect 9956 14016 10008 14068
rect 9128 13948 9180 14000
rect 11060 14016 11112 14068
rect 14004 14016 14056 14068
rect 10508 13948 10560 14000
rect 5816 13923 5868 13932
rect 2412 13744 2464 13796
rect 1492 13676 1544 13728
rect 2228 13676 2280 13728
rect 2964 13812 3016 13864
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 5816 13880 5868 13889
rect 6460 13880 6512 13932
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 7196 13880 7248 13932
rect 9404 13880 9456 13932
rect 10232 13880 10284 13932
rect 12072 13948 12124 14000
rect 12716 13923 12768 13932
rect 9496 13812 9548 13864
rect 2872 13719 2924 13728
rect 2872 13685 2902 13719
rect 2902 13685 2924 13719
rect 2872 13676 2924 13685
rect 3976 13676 4028 13728
rect 7012 13744 7064 13796
rect 4712 13676 4764 13728
rect 7196 13676 7248 13728
rect 8668 13744 8720 13796
rect 9864 13812 9916 13864
rect 9956 13812 10008 13864
rect 10416 13812 10468 13864
rect 9772 13744 9824 13796
rect 11336 13812 11388 13864
rect 12716 13889 12725 13923
rect 12725 13889 12759 13923
rect 12759 13889 12768 13923
rect 12716 13880 12768 13889
rect 12900 13880 12952 13932
rect 13084 13880 13136 13932
rect 13912 13948 13964 14000
rect 14464 13948 14516 14000
rect 15200 13948 15252 14000
rect 12072 13812 12124 13864
rect 12808 13812 12860 13864
rect 14004 13812 14056 13864
rect 11704 13744 11756 13796
rect 14280 13744 14332 13796
rect 16304 13744 16356 13796
rect 8576 13676 8628 13728
rect 9864 13676 9916 13728
rect 10968 13676 11020 13728
rect 11428 13676 11480 13728
rect 12900 13676 12952 13728
rect 16120 13676 16172 13728
rect 2924 13574 2976 13626
rect 2988 13574 3040 13626
rect 3052 13574 3104 13626
rect 3116 13574 3168 13626
rect 3180 13574 3232 13626
rect 6872 13574 6924 13626
rect 6936 13574 6988 13626
rect 7000 13574 7052 13626
rect 7064 13574 7116 13626
rect 7128 13574 7180 13626
rect 10820 13574 10872 13626
rect 10884 13574 10936 13626
rect 10948 13574 11000 13626
rect 11012 13574 11064 13626
rect 11076 13574 11128 13626
rect 14768 13574 14820 13626
rect 14832 13574 14884 13626
rect 14896 13574 14948 13626
rect 14960 13574 15012 13626
rect 15024 13574 15076 13626
rect 1860 13472 1912 13524
rect 2872 13404 2924 13456
rect 3700 13404 3752 13456
rect 5632 13472 5684 13524
rect 7012 13472 7064 13524
rect 7288 13472 7340 13524
rect 7564 13472 7616 13524
rect 7840 13472 7892 13524
rect 8484 13472 8536 13524
rect 9864 13472 9916 13524
rect 9956 13472 10008 13524
rect 11336 13472 11388 13524
rect 12164 13472 12216 13524
rect 1860 13336 1912 13388
rect 2228 13336 2280 13388
rect 3240 13336 3292 13388
rect 1492 13311 1544 13320
rect 1492 13277 1501 13311
rect 1501 13277 1535 13311
rect 1535 13277 1544 13311
rect 1492 13268 1544 13277
rect 3056 13268 3108 13320
rect 4528 13336 4580 13388
rect 5540 13336 5592 13388
rect 2044 13200 2096 13252
rect 3240 13200 3292 13252
rect 5448 13268 5500 13320
rect 5632 13268 5684 13320
rect 7288 13336 7340 13388
rect 7840 13336 7892 13388
rect 6736 13268 6788 13320
rect 7472 13268 7524 13320
rect 8208 13200 8260 13252
rect 9956 13336 10008 13388
rect 10416 13336 10468 13388
rect 12532 13404 12584 13456
rect 12716 13404 12768 13456
rect 12900 13515 12952 13524
rect 12900 13481 12909 13515
rect 12909 13481 12943 13515
rect 12943 13481 12952 13515
rect 12900 13472 12952 13481
rect 13176 13472 13228 13524
rect 14556 13472 14608 13524
rect 14740 13472 14792 13524
rect 15200 13472 15252 13524
rect 15384 13472 15436 13524
rect 8668 13268 8720 13320
rect 8760 13268 8812 13320
rect 10876 13268 10928 13320
rect 11152 13268 11204 13320
rect 11612 13268 11664 13320
rect 12440 13336 12492 13388
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 8484 13200 8536 13252
rect 8944 13200 8996 13252
rect 9036 13200 9088 13252
rect 10784 13200 10836 13252
rect 3056 13132 3108 13184
rect 5448 13132 5500 13184
rect 5908 13132 5960 13184
rect 6368 13132 6420 13184
rect 7104 13132 7156 13184
rect 9864 13132 9916 13184
rect 10416 13132 10468 13184
rect 10968 13132 11020 13184
rect 11796 13243 11848 13252
rect 11796 13209 11805 13243
rect 11805 13209 11839 13243
rect 11839 13209 11848 13243
rect 11796 13200 11848 13209
rect 12808 13200 12860 13252
rect 12992 13336 13044 13388
rect 13452 13268 13504 13320
rect 14556 13311 14608 13320
rect 14556 13277 14565 13311
rect 14565 13277 14599 13311
rect 14599 13277 14608 13311
rect 14556 13268 14608 13277
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 16028 13268 16080 13320
rect 12072 13132 12124 13184
rect 13544 13200 13596 13252
rect 13728 13132 13780 13184
rect 14188 13132 14240 13184
rect 16396 13132 16448 13184
rect 4898 13030 4950 13082
rect 4962 13030 5014 13082
rect 5026 13030 5078 13082
rect 5090 13030 5142 13082
rect 5154 13030 5206 13082
rect 8846 13030 8898 13082
rect 8910 13030 8962 13082
rect 8974 13030 9026 13082
rect 9038 13030 9090 13082
rect 9102 13030 9154 13082
rect 12794 13030 12846 13082
rect 12858 13030 12910 13082
rect 12922 13030 12974 13082
rect 12986 13030 13038 13082
rect 13050 13030 13102 13082
rect 480 12928 532 12980
rect 1124 12928 1176 12980
rect 2136 12928 2188 12980
rect 3056 12928 3108 12980
rect 2320 12860 2372 12912
rect 2044 12835 2096 12844
rect 2044 12801 2053 12835
rect 2053 12801 2087 12835
rect 2087 12801 2096 12835
rect 2044 12792 2096 12801
rect 2688 12792 2740 12844
rect 4160 12928 4212 12980
rect 4712 12928 4764 12980
rect 4896 12928 4948 12980
rect 5356 12928 5408 12980
rect 5908 12928 5960 12980
rect 7288 12928 7340 12980
rect 7840 12928 7892 12980
rect 9036 12928 9088 12980
rect 9128 12928 9180 12980
rect 5080 12860 5132 12912
rect 5448 12903 5500 12912
rect 5448 12869 5457 12903
rect 5457 12869 5491 12903
rect 5491 12869 5500 12903
rect 5448 12860 5500 12869
rect 6184 12860 6236 12912
rect 5172 12792 5224 12844
rect 5816 12792 5868 12844
rect 2228 12724 2280 12776
rect 3056 12724 3108 12776
rect 3240 12724 3292 12776
rect 4068 12724 4120 12776
rect 4528 12724 4580 12776
rect 2504 12656 2556 12708
rect 1952 12588 2004 12640
rect 2136 12588 2188 12640
rect 5356 12656 5408 12708
rect 5540 12656 5592 12708
rect 6000 12656 6052 12708
rect 4528 12588 4580 12640
rect 7564 12860 7616 12912
rect 8484 12860 8536 12912
rect 9772 12860 9824 12912
rect 9864 12860 9916 12912
rect 12256 12928 12308 12980
rect 12808 12928 12860 12980
rect 7748 12792 7800 12844
rect 7840 12835 7892 12844
rect 7840 12801 7849 12835
rect 7849 12801 7883 12835
rect 7883 12801 7892 12835
rect 7840 12792 7892 12801
rect 8852 12792 8904 12844
rect 9956 12792 10008 12844
rect 10324 12792 10376 12844
rect 10600 12792 10652 12844
rect 10692 12792 10744 12844
rect 10968 12835 11020 12844
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 11336 12792 11388 12844
rect 7104 12724 7156 12776
rect 7472 12724 7524 12776
rect 6368 12656 6420 12708
rect 9220 12724 9272 12776
rect 9496 12724 9548 12776
rect 7840 12656 7892 12708
rect 6552 12588 6604 12640
rect 8852 12588 8904 12640
rect 9312 12656 9364 12708
rect 10876 12724 10928 12776
rect 12532 12792 12584 12844
rect 12808 12792 12860 12844
rect 12992 12860 13044 12912
rect 13452 12860 13504 12912
rect 15200 12928 15252 12980
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 15660 12928 15712 12980
rect 14004 12860 14056 12912
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 14648 12792 14700 12844
rect 14832 12792 14884 12844
rect 15384 12792 15436 12844
rect 9496 12588 9548 12640
rect 10324 12588 10376 12640
rect 11796 12656 11848 12708
rect 12532 12656 12584 12708
rect 12992 12656 13044 12708
rect 12440 12588 12492 12640
rect 16304 12724 16356 12776
rect 14004 12656 14056 12708
rect 13360 12588 13412 12640
rect 13820 12588 13872 12640
rect 14096 12588 14148 12640
rect 14464 12588 14516 12640
rect 14740 12588 14792 12640
rect 15200 12588 15252 12640
rect 15752 12588 15804 12640
rect 2924 12486 2976 12538
rect 2988 12486 3040 12538
rect 3052 12486 3104 12538
rect 3116 12486 3168 12538
rect 3180 12486 3232 12538
rect 6872 12486 6924 12538
rect 6936 12486 6988 12538
rect 7000 12486 7052 12538
rect 7064 12486 7116 12538
rect 7128 12486 7180 12538
rect 10820 12486 10872 12538
rect 10884 12486 10936 12538
rect 10948 12486 11000 12538
rect 11012 12486 11064 12538
rect 11076 12486 11128 12538
rect 14768 12486 14820 12538
rect 14832 12486 14884 12538
rect 14896 12486 14948 12538
rect 14960 12486 15012 12538
rect 15024 12486 15076 12538
rect 2044 12384 2096 12436
rect 4160 12384 4212 12436
rect 296 12316 348 12368
rect 940 12248 992 12300
rect 3056 12316 3108 12368
rect 3424 12316 3476 12368
rect 3608 12316 3660 12368
rect 8668 12384 8720 12436
rect 9312 12384 9364 12436
rect 11336 12384 11388 12436
rect 2136 12248 2188 12300
rect 3148 12248 3200 12300
rect 3884 12248 3936 12300
rect 4436 12291 4488 12300
rect 4436 12257 4445 12291
rect 4445 12257 4479 12291
rect 4479 12257 4488 12291
rect 4436 12248 4488 12257
rect 7012 12316 7064 12368
rect 9680 12316 9732 12368
rect 13176 12384 13228 12436
rect 14004 12384 14056 12436
rect 14096 12384 14148 12436
rect 4988 12291 5040 12300
rect 4988 12257 4997 12291
rect 4997 12257 5031 12291
rect 5031 12257 5040 12291
rect 4988 12248 5040 12257
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 2596 12223 2648 12232
rect 2320 12180 2372 12189
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 3424 12180 3476 12232
rect 4804 12223 4856 12232
rect 4804 12189 4838 12223
rect 4838 12189 4856 12223
rect 4804 12180 4856 12189
rect 3884 12112 3936 12164
rect 6736 12248 6788 12300
rect 6920 12180 6972 12232
rect 8024 12180 8076 12232
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 10876 12248 10928 12300
rect 13084 12316 13136 12368
rect 13452 12316 13504 12368
rect 14648 12316 14700 12368
rect 15108 12384 15160 12436
rect 15384 12384 15436 12436
rect 15660 12316 15712 12368
rect 7012 12112 7064 12164
rect 8116 12112 8168 12164
rect 2688 12044 2740 12096
rect 5908 12044 5960 12096
rect 6276 12044 6328 12096
rect 6828 12044 6880 12096
rect 7196 12044 7248 12096
rect 8208 12044 8260 12096
rect 8484 12044 8536 12096
rect 9956 12155 10008 12164
rect 9956 12121 9990 12155
rect 9990 12121 10008 12155
rect 13636 12180 13688 12232
rect 13912 12248 13964 12300
rect 14096 12248 14148 12300
rect 14372 12248 14424 12300
rect 9956 12112 10008 12121
rect 14648 12180 14700 12232
rect 15108 12180 15160 12232
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15936 12223 15988 12232
rect 15476 12180 15528 12189
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 14924 12112 14976 12164
rect 11060 12087 11112 12096
rect 11060 12053 11069 12087
rect 11069 12053 11103 12087
rect 11103 12053 11112 12087
rect 11060 12044 11112 12053
rect 11152 12044 11204 12096
rect 12900 12044 12952 12096
rect 13268 12044 13320 12096
rect 15568 12112 15620 12164
rect 15936 12044 15988 12096
rect 16396 12044 16448 12096
rect 4898 11942 4950 11994
rect 4962 11942 5014 11994
rect 5026 11942 5078 11994
rect 5090 11942 5142 11994
rect 5154 11942 5206 11994
rect 8846 11942 8898 11994
rect 8910 11942 8962 11994
rect 8974 11942 9026 11994
rect 9038 11942 9090 11994
rect 9102 11942 9154 11994
rect 12794 11942 12846 11994
rect 12858 11942 12910 11994
rect 12922 11942 12974 11994
rect 12986 11942 13038 11994
rect 13050 11942 13102 11994
rect 2780 11840 2832 11892
rect 2964 11840 3016 11892
rect 3424 11840 3476 11892
rect 4712 11883 4764 11892
rect 4712 11849 4721 11883
rect 4721 11849 4755 11883
rect 4755 11849 4764 11883
rect 4712 11840 4764 11849
rect 5080 11840 5132 11892
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 2136 11704 2188 11756
rect 3240 11704 3292 11756
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 5172 11747 5224 11756
rect 5172 11713 5181 11747
rect 5181 11713 5215 11747
rect 5215 11713 5224 11747
rect 5172 11704 5224 11713
rect 2228 11636 2280 11688
rect 3056 11568 3108 11620
rect 3516 11611 3568 11620
rect 3516 11577 3525 11611
rect 3525 11577 3559 11611
rect 3559 11577 3568 11611
rect 3516 11568 3568 11577
rect 388 11500 440 11552
rect 2044 11500 2096 11552
rect 2320 11500 2372 11552
rect 5172 11500 5224 11552
rect 5724 11704 5776 11756
rect 6460 11704 6512 11756
rect 8116 11772 8168 11824
rect 8208 11704 8260 11756
rect 9588 11840 9640 11892
rect 10324 11840 10376 11892
rect 10508 11840 10560 11892
rect 10600 11883 10652 11892
rect 10600 11849 10609 11883
rect 10609 11849 10643 11883
rect 10643 11849 10652 11883
rect 10600 11840 10652 11849
rect 10784 11840 10836 11892
rect 11336 11840 11388 11892
rect 11428 11840 11480 11892
rect 13268 11840 13320 11892
rect 13728 11840 13780 11892
rect 13176 11772 13228 11824
rect 13452 11772 13504 11824
rect 5816 11679 5868 11688
rect 5816 11645 5825 11679
rect 5825 11645 5859 11679
rect 5859 11645 5868 11679
rect 5816 11636 5868 11645
rect 9128 11704 9180 11756
rect 11612 11704 11664 11756
rect 12072 11704 12124 11756
rect 6276 11568 6328 11620
rect 8392 11568 8444 11620
rect 12716 11704 12768 11756
rect 15292 11840 15344 11892
rect 14372 11772 14424 11824
rect 14740 11815 14792 11824
rect 14740 11781 14749 11815
rect 14749 11781 14783 11815
rect 14783 11781 14792 11815
rect 14740 11772 14792 11781
rect 15292 11704 15344 11756
rect 5632 11500 5684 11552
rect 7472 11500 7524 11552
rect 10232 11500 10284 11552
rect 14096 11636 14148 11688
rect 14648 11636 14700 11688
rect 13268 11568 13320 11620
rect 13820 11500 13872 11552
rect 14188 11500 14240 11552
rect 16120 11500 16172 11552
rect 2924 11398 2976 11450
rect 2988 11398 3040 11450
rect 3052 11398 3104 11450
rect 3116 11398 3168 11450
rect 3180 11398 3232 11450
rect 6872 11398 6924 11450
rect 6936 11398 6988 11450
rect 7000 11398 7052 11450
rect 7064 11398 7116 11450
rect 7128 11398 7180 11450
rect 10820 11398 10872 11450
rect 10884 11398 10936 11450
rect 10948 11398 11000 11450
rect 11012 11398 11064 11450
rect 11076 11398 11128 11450
rect 14768 11398 14820 11450
rect 14832 11398 14884 11450
rect 14896 11398 14948 11450
rect 14960 11398 15012 11450
rect 15024 11398 15076 11450
rect 2964 11160 3016 11212
rect 10784 11296 10836 11348
rect 4068 11228 4120 11280
rect 4252 11160 4304 11212
rect 5908 11228 5960 11280
rect 6276 11228 6328 11280
rect 6460 11228 6512 11280
rect 7472 11228 7524 11280
rect 10140 11228 10192 11280
rect 10324 11228 10376 11280
rect 10416 11228 10468 11280
rect 10600 11228 10652 11280
rect 7380 11160 7432 11212
rect 7840 11160 7892 11212
rect 8668 11160 8720 11212
rect 7104 11092 7156 11144
rect 1860 11024 1912 11076
rect 3424 11024 3476 11076
rect 4160 11024 4212 11076
rect 6460 11024 6512 11076
rect 7840 11024 7892 11076
rect 9956 11092 10008 11144
rect 10692 11092 10744 11144
rect 11520 11092 11572 11144
rect 9036 11024 9088 11076
rect 9588 11024 9640 11076
rect 9680 11024 9732 11076
rect 10876 11024 10928 11076
rect 11244 11024 11296 11076
rect 11428 11024 11480 11076
rect 11980 11296 12032 11348
rect 12164 11339 12216 11348
rect 12164 11305 12173 11339
rect 12173 11305 12207 11339
rect 12207 11305 12216 11339
rect 12164 11296 12216 11305
rect 12624 11296 12676 11348
rect 12808 11296 12860 11348
rect 13176 11228 13228 11280
rect 14096 11296 14148 11348
rect 15200 11296 15252 11348
rect 16120 11296 16172 11348
rect 16856 11296 16908 11348
rect 12072 11092 12124 11144
rect 12164 11092 12216 11144
rect 12808 11092 12860 11144
rect 13084 11092 13136 11144
rect 13636 11160 13688 11212
rect 14924 11228 14976 11280
rect 13728 11092 13780 11144
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 14648 11092 14700 11144
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 16856 11160 16908 11212
rect 1584 10956 1636 11008
rect 2596 10956 2648 11008
rect 3332 10956 3384 11008
rect 5540 10956 5592 11008
rect 7288 10956 7340 11008
rect 9128 10956 9180 11008
rect 9772 10956 9824 11008
rect 10600 10956 10652 11008
rect 12992 10956 13044 11008
rect 13360 10956 13412 11008
rect 14556 11024 14608 11076
rect 14188 10956 14240 11008
rect 4898 10854 4950 10906
rect 4962 10854 5014 10906
rect 5026 10854 5078 10906
rect 5090 10854 5142 10906
rect 5154 10854 5206 10906
rect 8846 10854 8898 10906
rect 8910 10854 8962 10906
rect 8974 10854 9026 10906
rect 9038 10854 9090 10906
rect 9102 10854 9154 10906
rect 12794 10854 12846 10906
rect 12858 10854 12910 10906
rect 12922 10854 12974 10906
rect 12986 10854 13038 10906
rect 13050 10854 13102 10906
rect 1768 10795 1820 10804
rect 1768 10761 1777 10795
rect 1777 10761 1811 10795
rect 1811 10761 1820 10795
rect 1768 10752 1820 10761
rect 2136 10752 2188 10804
rect 4620 10752 4672 10804
rect 10968 10752 11020 10804
rect 12532 10752 12584 10804
rect 13176 10752 13228 10804
rect 14188 10752 14240 10804
rect 13728 10727 13780 10736
rect 13728 10693 13737 10727
rect 13737 10693 13771 10727
rect 13771 10693 13780 10727
rect 13728 10684 13780 10693
rect 1768 10616 1820 10668
rect 1584 10548 1636 10600
rect 2688 10548 2740 10600
rect 2872 10659 2924 10668
rect 2872 10625 2881 10659
rect 2881 10625 2915 10659
rect 2915 10625 2924 10659
rect 2872 10616 2924 10625
rect 3700 10616 3752 10668
rect 5172 10548 5224 10600
rect 5356 10591 5408 10600
rect 5356 10557 5365 10591
rect 5365 10557 5399 10591
rect 5399 10557 5408 10591
rect 5356 10548 5408 10557
rect 8484 10616 8536 10668
rect 8760 10616 8812 10668
rect 9956 10616 10008 10668
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10140 10616 10192 10625
rect 11152 10616 11204 10668
rect 12808 10616 12860 10668
rect 13636 10659 13688 10668
rect 13636 10625 13644 10659
rect 13644 10625 13678 10659
rect 13678 10625 13688 10659
rect 13636 10616 13688 10625
rect 940 10412 992 10464
rect 5080 10480 5132 10532
rect 5540 10480 5592 10532
rect 6184 10480 6236 10532
rect 10600 10548 10652 10600
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 12532 10548 12584 10600
rect 14096 10616 14148 10668
rect 14556 10684 14608 10736
rect 14740 10727 14792 10736
rect 14740 10693 14749 10727
rect 14749 10693 14783 10727
rect 14783 10693 14792 10727
rect 15292 10752 15344 10804
rect 16120 10752 16172 10804
rect 14740 10684 14792 10693
rect 14832 10659 14884 10668
rect 14832 10625 14841 10659
rect 14841 10625 14875 10659
rect 14875 10625 14884 10659
rect 14832 10616 14884 10625
rect 7932 10480 7984 10532
rect 4896 10412 4948 10464
rect 11244 10480 11296 10532
rect 13452 10480 13504 10532
rect 14648 10548 14700 10600
rect 15108 10616 15160 10668
rect 15016 10548 15068 10600
rect 15476 10523 15528 10532
rect 15476 10489 15485 10523
rect 15485 10489 15519 10523
rect 15519 10489 15528 10523
rect 15476 10480 15528 10489
rect 15660 10480 15712 10532
rect 8392 10412 8444 10464
rect 8576 10412 8628 10464
rect 10140 10412 10192 10464
rect 10508 10412 10560 10464
rect 10784 10412 10836 10464
rect 12256 10412 12308 10464
rect 12440 10412 12492 10464
rect 13176 10412 13228 10464
rect 13544 10412 13596 10464
rect 14096 10412 14148 10464
rect 14188 10412 14240 10464
rect 16856 10412 16908 10464
rect 2924 10310 2976 10362
rect 2988 10310 3040 10362
rect 3052 10310 3104 10362
rect 3116 10310 3168 10362
rect 3180 10310 3232 10362
rect 6872 10310 6924 10362
rect 6936 10310 6988 10362
rect 7000 10310 7052 10362
rect 7064 10310 7116 10362
rect 7128 10310 7180 10362
rect 10820 10310 10872 10362
rect 10884 10310 10936 10362
rect 10948 10310 11000 10362
rect 11012 10310 11064 10362
rect 11076 10310 11128 10362
rect 14768 10310 14820 10362
rect 14832 10310 14884 10362
rect 14896 10310 14948 10362
rect 14960 10310 15012 10362
rect 15024 10310 15076 10362
rect 3884 10251 3936 10260
rect 3884 10217 3893 10251
rect 3893 10217 3927 10251
rect 3927 10217 3936 10251
rect 3884 10208 3936 10217
rect 1400 10140 1452 10192
rect 5172 10208 5224 10260
rect 8116 10251 8168 10260
rect 8116 10217 8125 10251
rect 8125 10217 8159 10251
rect 8159 10217 8168 10251
rect 8116 10208 8168 10217
rect 9312 10208 9364 10260
rect 11336 10208 11388 10260
rect 11520 10208 11572 10260
rect 11980 10208 12032 10260
rect 1492 10115 1544 10124
rect 1492 10081 1501 10115
rect 1501 10081 1535 10115
rect 1535 10081 1544 10115
rect 1492 10072 1544 10081
rect 3148 10072 3200 10124
rect 5724 10140 5776 10192
rect 5908 10140 5960 10192
rect 6184 10140 6236 10192
rect 8300 10140 8352 10192
rect 9956 10140 10008 10192
rect 12808 10208 12860 10260
rect 13912 10208 13964 10260
rect 4068 10072 4120 10124
rect 5080 10072 5132 10124
rect 9036 10072 9088 10124
rect 14096 10140 14148 10192
rect 14556 10140 14608 10192
rect 14740 10208 14792 10260
rect 15476 10208 15528 10260
rect 15660 10208 15712 10260
rect 16396 10208 16448 10260
rect 3700 10004 3752 10056
rect 2780 9936 2832 9988
rect 3332 9936 3384 9988
rect 4252 10004 4304 10056
rect 6736 10004 6788 10056
rect 7196 10004 7248 10056
rect 7932 10004 7984 10056
rect 8760 10004 8812 10056
rect 11428 10004 11480 10056
rect 12072 10004 12124 10056
rect 13268 10072 13320 10124
rect 12532 10004 12584 10056
rect 12808 10004 12860 10056
rect 12992 10047 13044 10056
rect 12992 10013 13001 10047
rect 13001 10013 13035 10047
rect 13035 10013 13044 10047
rect 12992 10004 13044 10013
rect 14556 10047 14608 10056
rect 6092 9936 6144 9988
rect 10508 9936 10560 9988
rect 4160 9868 4212 9920
rect 6368 9868 6420 9920
rect 8576 9868 8628 9920
rect 13636 9936 13688 9988
rect 13820 9936 13872 9988
rect 14556 10013 14565 10047
rect 14565 10013 14599 10047
rect 14599 10013 14608 10047
rect 14556 10004 14608 10013
rect 15476 10072 15528 10124
rect 16212 10072 16264 10124
rect 14924 10047 14976 10056
rect 14924 10013 14947 10047
rect 14947 10013 14976 10047
rect 14924 10004 14976 10013
rect 16856 10004 16908 10056
rect 15752 9936 15804 9988
rect 16396 9936 16448 9988
rect 11428 9868 11480 9920
rect 14280 9868 14332 9920
rect 14372 9911 14424 9920
rect 14372 9877 14381 9911
rect 14381 9877 14415 9911
rect 14415 9877 14424 9911
rect 14372 9868 14424 9877
rect 14556 9868 14608 9920
rect 4898 9766 4950 9818
rect 4962 9766 5014 9818
rect 5026 9766 5078 9818
rect 5090 9766 5142 9818
rect 5154 9766 5206 9818
rect 8846 9766 8898 9818
rect 8910 9766 8962 9818
rect 8974 9766 9026 9818
rect 9038 9766 9090 9818
rect 9102 9766 9154 9818
rect 12794 9766 12846 9818
rect 12858 9766 12910 9818
rect 12922 9766 12974 9818
rect 12986 9766 13038 9818
rect 13050 9766 13102 9818
rect 1032 9664 1084 9716
rect 1584 9664 1636 9716
rect 4068 9664 4120 9716
rect 9588 9664 9640 9716
rect 10324 9664 10376 9716
rect 10600 9664 10652 9716
rect 11336 9664 11388 9716
rect 2320 9596 2372 9648
rect 3240 9528 3292 9580
rect 5908 9596 5960 9648
rect 2136 9460 2188 9512
rect 3148 9460 3200 9512
rect 2780 9392 2832 9444
rect 3884 9460 3936 9512
rect 5448 9528 5500 9580
rect 7288 9596 7340 9648
rect 8116 9596 8168 9648
rect 8852 9596 8904 9648
rect 11980 9596 12032 9648
rect 6092 9460 6144 9512
rect 6368 9460 6420 9512
rect 11244 9528 11296 9580
rect 11612 9528 11664 9580
rect 12348 9528 12400 9580
rect 13268 9664 13320 9716
rect 12900 9596 12952 9648
rect 14832 9664 14884 9716
rect 15292 9664 15344 9716
rect 15936 9664 15988 9716
rect 15200 9528 15252 9580
rect 9956 9460 10008 9512
rect 10984 9460 11036 9512
rect 11336 9460 11388 9512
rect 13360 9503 13412 9512
rect 13360 9469 13369 9503
rect 13369 9469 13403 9503
rect 13403 9469 13412 9503
rect 13360 9460 13412 9469
rect 9404 9392 9456 9444
rect 11520 9392 11572 9444
rect 12532 9392 12584 9444
rect 12900 9435 12952 9444
rect 12900 9401 12909 9435
rect 12909 9401 12943 9435
rect 12943 9401 12952 9435
rect 12900 9392 12952 9401
rect 15660 9571 15712 9580
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 15660 9528 15712 9537
rect 4160 9324 4212 9376
rect 4804 9324 4856 9376
rect 5448 9324 5500 9376
rect 6828 9324 6880 9376
rect 8668 9324 8720 9376
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 10600 9324 10652 9376
rect 15660 9324 15712 9376
rect 2924 9222 2976 9274
rect 2988 9222 3040 9274
rect 3052 9222 3104 9274
rect 3116 9222 3168 9274
rect 3180 9222 3232 9274
rect 6872 9222 6924 9274
rect 6936 9222 6988 9274
rect 7000 9222 7052 9274
rect 7064 9222 7116 9274
rect 7128 9222 7180 9274
rect 10820 9222 10872 9274
rect 10884 9222 10936 9274
rect 10948 9222 11000 9274
rect 11012 9222 11064 9274
rect 11076 9222 11128 9274
rect 14768 9222 14820 9274
rect 14832 9222 14884 9274
rect 14896 9222 14948 9274
rect 14960 9222 15012 9274
rect 15024 9222 15076 9274
rect 6092 9120 6144 9172
rect 6276 9163 6328 9172
rect 6276 9129 6285 9163
rect 6285 9129 6319 9163
rect 6319 9129 6328 9163
rect 6276 9120 6328 9129
rect 7932 9120 7984 9172
rect 8576 9120 8628 9172
rect 2136 8984 2188 9036
rect 9220 9052 9272 9104
rect 10600 9052 10652 9104
rect 4436 8984 4488 9036
rect 5816 8984 5868 9036
rect 6552 8984 6604 9036
rect 8852 8984 8904 9036
rect 6736 8916 6788 8968
rect 7104 8916 7156 8968
rect 1032 8848 1084 8900
rect 3884 8848 3936 8900
rect 6644 8848 6696 8900
rect 7472 8848 7524 8900
rect 7748 8916 7800 8968
rect 9588 8984 9640 9036
rect 11336 9052 11388 9104
rect 12532 9052 12584 9104
rect 12808 9052 12860 9104
rect 11152 8984 11204 9036
rect 12716 8984 12768 9036
rect 12992 8916 13044 8968
rect 14096 8984 14148 9036
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 15568 9120 15620 9172
rect 15936 9052 15988 9104
rect 14832 8984 14884 9036
rect 13728 8916 13780 8968
rect 14004 8916 14056 8968
rect 14648 8916 14700 8968
rect 15016 8916 15068 8968
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 6092 8780 6144 8832
rect 9312 8780 9364 8832
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 10784 8780 10836 8789
rect 11152 8848 11204 8900
rect 11428 8848 11480 8900
rect 11980 8848 12032 8900
rect 12348 8848 12400 8900
rect 15752 8916 15804 8968
rect 16212 8916 16264 8968
rect 15384 8780 15436 8832
rect 4898 8678 4950 8730
rect 4962 8678 5014 8730
rect 5026 8678 5078 8730
rect 5090 8678 5142 8730
rect 5154 8678 5206 8730
rect 8846 8678 8898 8730
rect 8910 8678 8962 8730
rect 8974 8678 9026 8730
rect 9038 8678 9090 8730
rect 9102 8678 9154 8730
rect 12794 8678 12846 8730
rect 12858 8678 12910 8730
rect 12922 8678 12974 8730
rect 12986 8678 13038 8730
rect 13050 8678 13102 8730
rect 3608 8576 3660 8628
rect 9588 8576 9640 8628
rect 5448 8508 5500 8560
rect 6368 8508 6420 8560
rect 12440 8576 12492 8628
rect 13452 8576 13504 8628
rect 13544 8576 13596 8628
rect 14740 8576 14792 8628
rect 10876 8508 10928 8560
rect 12900 8508 12952 8560
rect 3608 8440 3660 8492
rect 5172 8440 5224 8492
rect 8300 8440 8352 8492
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 4068 8415 4120 8424
rect 2044 8236 2096 8288
rect 2320 8236 2372 8288
rect 4068 8381 4077 8415
rect 4077 8381 4111 8415
rect 4111 8381 4120 8415
rect 4068 8372 4120 8381
rect 4436 8372 4488 8424
rect 6368 8415 6420 8424
rect 6368 8381 6377 8415
rect 6377 8381 6411 8415
rect 6411 8381 6420 8415
rect 6368 8372 6420 8381
rect 5080 8304 5132 8356
rect 9588 8372 9640 8424
rect 12348 8440 12400 8492
rect 12808 8440 12860 8492
rect 13728 8551 13780 8560
rect 13728 8517 13737 8551
rect 13737 8517 13771 8551
rect 13771 8517 13780 8551
rect 13728 8508 13780 8517
rect 14648 8508 14700 8560
rect 11336 8372 11388 8424
rect 6092 8236 6144 8288
rect 8300 8236 8352 8288
rect 11336 8236 11388 8288
rect 11520 8236 11572 8288
rect 14096 8372 14148 8424
rect 13084 8304 13136 8356
rect 13544 8304 13596 8356
rect 13636 8304 13688 8356
rect 14740 8372 14792 8424
rect 16396 8440 16448 8492
rect 15752 8372 15804 8424
rect 15108 8304 15160 8356
rect 15292 8304 15344 8356
rect 15016 8236 15068 8288
rect 17684 8236 17736 8288
rect 2924 8134 2976 8186
rect 2988 8134 3040 8186
rect 3052 8134 3104 8186
rect 3116 8134 3168 8186
rect 3180 8134 3232 8186
rect 6872 8134 6924 8186
rect 6936 8134 6988 8186
rect 7000 8134 7052 8186
rect 7064 8134 7116 8186
rect 7128 8134 7180 8186
rect 10820 8134 10872 8186
rect 10884 8134 10936 8186
rect 10948 8134 11000 8186
rect 11012 8134 11064 8186
rect 11076 8134 11128 8186
rect 14768 8134 14820 8186
rect 14832 8134 14884 8186
rect 14896 8134 14948 8186
rect 14960 8134 15012 8186
rect 15024 8134 15076 8186
rect 1952 8032 2004 8084
rect 2320 8032 2372 8084
rect 4068 8032 4120 8084
rect 6184 8032 6236 8084
rect 7840 8032 7892 8084
rect 4436 7964 4488 8016
rect 10784 8032 10836 8084
rect 11980 8032 12032 8084
rect 5080 7828 5132 7880
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 7564 7828 7616 7880
rect 8024 7828 8076 7880
rect 4804 7760 4856 7812
rect 8392 7760 8444 7812
rect 9404 7896 9456 7948
rect 9772 7896 9824 7948
rect 13360 7964 13412 8016
rect 13544 7964 13596 8016
rect 11336 7896 11388 7948
rect 12348 7896 12400 7948
rect 9220 7828 9272 7880
rect 9312 7828 9364 7880
rect 10416 7803 10468 7812
rect 2504 7692 2556 7744
rect 3332 7692 3384 7744
rect 4160 7692 4212 7744
rect 4620 7692 4672 7744
rect 5356 7692 5408 7744
rect 7288 7692 7340 7744
rect 7932 7692 7984 7744
rect 8668 7692 8720 7744
rect 9036 7692 9088 7744
rect 9864 7692 9916 7744
rect 10416 7769 10425 7803
rect 10425 7769 10459 7803
rect 10459 7769 10468 7803
rect 10416 7760 10468 7769
rect 10600 7760 10652 7812
rect 10784 7760 10836 7812
rect 13452 7828 13504 7880
rect 13728 7760 13780 7812
rect 13912 7896 13964 7948
rect 14740 7828 14792 7880
rect 15384 7828 15436 7880
rect 16212 7828 16264 7880
rect 16672 7760 16724 7812
rect 11336 7692 11388 7744
rect 11520 7692 11572 7744
rect 11980 7692 12032 7744
rect 13912 7692 13964 7744
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 14832 7692 14884 7744
rect 16396 7692 16448 7744
rect 4898 7590 4950 7642
rect 4962 7590 5014 7642
rect 5026 7590 5078 7642
rect 5090 7590 5142 7642
rect 5154 7590 5206 7642
rect 8846 7590 8898 7642
rect 8910 7590 8962 7642
rect 8974 7590 9026 7642
rect 9038 7590 9090 7642
rect 9102 7590 9154 7642
rect 12794 7590 12846 7642
rect 12858 7590 12910 7642
rect 12922 7590 12974 7642
rect 12986 7590 13038 7642
rect 13050 7590 13102 7642
rect 1952 7488 2004 7540
rect 9496 7488 9548 7540
rect 1492 7352 1544 7404
rect 7380 7420 7432 7472
rect 7840 7463 7892 7472
rect 7840 7429 7849 7463
rect 7849 7429 7883 7463
rect 7883 7429 7892 7463
rect 7840 7420 7892 7429
rect 7932 7420 7984 7472
rect 11428 7488 11480 7540
rect 12072 7488 12124 7540
rect 12900 7488 12952 7540
rect 2688 7284 2740 7336
rect 6000 7352 6052 7404
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 7748 7352 7800 7404
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 5632 7284 5684 7336
rect 6276 7284 6328 7336
rect 7288 7284 7340 7336
rect 11980 7420 12032 7472
rect 12532 7420 12584 7472
rect 13912 7488 13964 7540
rect 15384 7488 15436 7540
rect 16948 7488 17000 7540
rect 11888 7352 11940 7404
rect 13360 7420 13412 7472
rect 14740 7420 14792 7472
rect 15016 7420 15068 7472
rect 12992 7352 13044 7404
rect 14832 7352 14884 7404
rect 11244 7284 11296 7336
rect 11980 7284 12032 7336
rect 7932 7216 7984 7268
rect 8944 7216 8996 7268
rect 9772 7216 9824 7268
rect 10692 7259 10744 7268
rect 10692 7225 10701 7259
rect 10701 7225 10735 7259
rect 10735 7225 10744 7259
rect 10692 7216 10744 7225
rect 11612 7216 11664 7268
rect 15384 7352 15436 7404
rect 12808 7216 12860 7268
rect 3700 7148 3752 7200
rect 4068 7148 4120 7200
rect 7472 7148 7524 7200
rect 8392 7148 8444 7200
rect 8576 7148 8628 7200
rect 9588 7148 9640 7200
rect 12716 7148 12768 7200
rect 13176 7148 13228 7200
rect 15568 7216 15620 7268
rect 15752 7216 15804 7268
rect 16212 7148 16264 7200
rect 2924 7046 2976 7098
rect 2988 7046 3040 7098
rect 3052 7046 3104 7098
rect 3116 7046 3168 7098
rect 3180 7046 3232 7098
rect 6872 7046 6924 7098
rect 6936 7046 6988 7098
rect 7000 7046 7052 7098
rect 7064 7046 7116 7098
rect 7128 7046 7180 7098
rect 10820 7046 10872 7098
rect 10884 7046 10936 7098
rect 10948 7046 11000 7098
rect 11012 7046 11064 7098
rect 11076 7046 11128 7098
rect 14768 7046 14820 7098
rect 14832 7046 14884 7098
rect 14896 7046 14948 7098
rect 14960 7046 15012 7098
rect 15024 7046 15076 7098
rect 2228 6944 2280 6996
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 1768 6808 1820 6860
rect 4344 6808 4396 6860
rect 7472 6944 7524 6996
rect 5172 6876 5224 6928
rect 7564 6876 7616 6928
rect 8760 6944 8812 6996
rect 9588 6944 9640 6996
rect 5172 6740 5224 6792
rect 5448 6740 5500 6792
rect 7840 6808 7892 6860
rect 8024 6783 8076 6792
rect 4804 6672 4856 6724
rect 4068 6604 4120 6656
rect 4620 6604 4672 6656
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 6460 6672 6512 6724
rect 8852 6808 8904 6860
rect 9404 6808 9456 6860
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 9312 6740 9364 6792
rect 11428 6944 11480 6996
rect 13268 6944 13320 6996
rect 14740 6944 14792 6996
rect 16304 6944 16356 6996
rect 12624 6876 12676 6928
rect 12532 6808 12584 6860
rect 15200 6876 15252 6928
rect 16672 6876 16724 6928
rect 10784 6740 10836 6792
rect 10876 6740 10928 6792
rect 11612 6740 11664 6792
rect 12256 6740 12308 6792
rect 12900 6740 12952 6792
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 14188 6740 14240 6792
rect 14740 6740 14792 6792
rect 15200 6740 15252 6792
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 9128 6672 9180 6724
rect 11428 6672 11480 6724
rect 6736 6604 6788 6656
rect 9588 6604 9640 6656
rect 10048 6604 10100 6656
rect 10692 6604 10744 6656
rect 10784 6604 10836 6656
rect 11980 6604 12032 6656
rect 12532 6604 12584 6656
rect 13452 6647 13504 6656
rect 13452 6613 13461 6647
rect 13461 6613 13495 6647
rect 13495 6613 13504 6647
rect 13452 6604 13504 6613
rect 13820 6604 13872 6656
rect 15568 6604 15620 6656
rect 4898 6502 4950 6554
rect 4962 6502 5014 6554
rect 5026 6502 5078 6554
rect 5090 6502 5142 6554
rect 5154 6502 5206 6554
rect 8846 6502 8898 6554
rect 8910 6502 8962 6554
rect 8974 6502 9026 6554
rect 9038 6502 9090 6554
rect 9102 6502 9154 6554
rect 12794 6502 12846 6554
rect 12858 6502 12910 6554
rect 12922 6502 12974 6554
rect 12986 6502 13038 6554
rect 13050 6502 13102 6554
rect 2780 6400 2832 6452
rect 7656 6400 7708 6452
rect 8760 6443 8812 6452
rect 8760 6409 8769 6443
rect 8769 6409 8803 6443
rect 8803 6409 8812 6443
rect 8760 6400 8812 6409
rect 4344 6332 4396 6384
rect 8208 6332 8260 6384
rect 1492 6264 1544 6316
rect 5908 6264 5960 6316
rect 6460 6264 6512 6316
rect 3700 6196 3752 6248
rect 5356 6196 5408 6248
rect 5540 6196 5592 6248
rect 5816 6196 5868 6248
rect 7104 6264 7156 6316
rect 7196 6264 7248 6316
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 10416 6400 10468 6452
rect 13084 6400 13136 6452
rect 11520 6332 11572 6384
rect 11980 6332 12032 6384
rect 9312 6264 9364 6316
rect 11152 6264 11204 6316
rect 8944 6196 8996 6248
rect 10324 6196 10376 6248
rect 13360 6264 13412 6316
rect 14648 6332 14700 6384
rect 11520 6239 11572 6248
rect 11520 6205 11529 6239
rect 11529 6205 11563 6239
rect 11563 6205 11572 6239
rect 11520 6196 11572 6205
rect 1492 6060 1544 6112
rect 3332 6103 3384 6112
rect 3332 6069 3341 6103
rect 3341 6069 3375 6103
rect 3375 6069 3384 6103
rect 7380 6128 7432 6180
rect 3332 6060 3384 6069
rect 5356 6060 5408 6112
rect 6552 6060 6604 6112
rect 10324 6060 10376 6112
rect 12716 6128 12768 6180
rect 12164 6060 12216 6112
rect 12532 6060 12584 6112
rect 13268 6060 13320 6112
rect 13544 6060 13596 6112
rect 14556 6264 14608 6316
rect 17500 6332 17552 6384
rect 17132 6264 17184 6316
rect 14096 6128 14148 6180
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 2924 5958 2976 6010
rect 2988 5958 3040 6010
rect 3052 5958 3104 6010
rect 3116 5958 3168 6010
rect 3180 5958 3232 6010
rect 6872 5958 6924 6010
rect 6936 5958 6988 6010
rect 7000 5958 7052 6010
rect 7064 5958 7116 6010
rect 7128 5958 7180 6010
rect 10820 5958 10872 6010
rect 10884 5958 10936 6010
rect 10948 5958 11000 6010
rect 11012 5958 11064 6010
rect 11076 5958 11128 6010
rect 14768 5958 14820 6010
rect 14832 5958 14884 6010
rect 14896 5958 14948 6010
rect 14960 5958 15012 6010
rect 15024 5958 15076 6010
rect 1492 5763 1544 5772
rect 1492 5729 1501 5763
rect 1501 5729 1535 5763
rect 1535 5729 1544 5763
rect 1492 5720 1544 5729
rect 6552 5856 6604 5908
rect 6736 5899 6788 5908
rect 6736 5865 6745 5899
rect 6745 5865 6779 5899
rect 6779 5865 6788 5899
rect 6736 5856 6788 5865
rect 7380 5856 7432 5908
rect 7840 5856 7892 5908
rect 7932 5856 7984 5908
rect 3332 5788 3384 5840
rect 8852 5788 8904 5840
rect 9680 5788 9732 5840
rect 3516 5720 3568 5772
rect 3332 5652 3384 5704
rect 4068 5652 4120 5704
rect 6644 5720 6696 5772
rect 5540 5652 5592 5704
rect 7932 5652 7984 5704
rect 8484 5720 8536 5772
rect 8116 5652 8168 5704
rect 9220 5652 9272 5704
rect 9772 5652 9824 5704
rect 2044 5516 2096 5568
rect 2780 5516 2832 5568
rect 3516 5516 3568 5568
rect 3700 5516 3752 5568
rect 4068 5516 4120 5568
rect 7656 5516 7708 5568
rect 8116 5516 8168 5568
rect 8484 5584 8536 5636
rect 9036 5516 9088 5568
rect 9312 5584 9364 5636
rect 9864 5516 9916 5568
rect 10232 5788 10284 5840
rect 10508 5788 10560 5840
rect 11888 5856 11940 5908
rect 12348 5856 12400 5908
rect 13452 5856 13504 5908
rect 14464 5899 14516 5908
rect 14464 5865 14473 5899
rect 14473 5865 14507 5899
rect 14507 5865 14516 5899
rect 14464 5856 14516 5865
rect 15108 5856 15160 5908
rect 10784 5720 10836 5772
rect 12440 5788 12492 5840
rect 12532 5788 12584 5840
rect 15384 5788 15436 5840
rect 11888 5720 11940 5772
rect 12624 5720 12676 5772
rect 13084 5720 13136 5772
rect 13544 5720 13596 5772
rect 13728 5720 13780 5772
rect 14556 5720 14608 5772
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 15844 5695 15896 5704
rect 11612 5584 11664 5636
rect 11428 5516 11480 5568
rect 12072 5516 12124 5568
rect 12808 5627 12860 5636
rect 12808 5593 12817 5627
rect 12817 5593 12851 5627
rect 12851 5593 12860 5627
rect 12808 5584 12860 5593
rect 12440 5516 12492 5568
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 13360 5516 13412 5568
rect 16028 5584 16080 5636
rect 4898 5414 4950 5466
rect 4962 5414 5014 5466
rect 5026 5414 5078 5466
rect 5090 5414 5142 5466
rect 5154 5414 5206 5466
rect 8846 5414 8898 5466
rect 8910 5414 8962 5466
rect 8974 5414 9026 5466
rect 9038 5414 9090 5466
rect 9102 5414 9154 5466
rect 12794 5414 12846 5466
rect 12858 5414 12910 5466
rect 12922 5414 12974 5466
rect 12986 5414 13038 5466
rect 13050 5414 13102 5466
rect 1952 5312 2004 5364
rect 2596 5312 2648 5364
rect 848 5244 900 5296
rect 6460 5312 6512 5364
rect 6552 5312 6604 5364
rect 7840 5312 7892 5364
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 1860 5176 1912 5228
rect 1768 5151 1820 5160
rect 1768 5117 1777 5151
rect 1777 5117 1811 5151
rect 1811 5117 1820 5151
rect 1768 5108 1820 5117
rect 5080 5176 5132 5228
rect 3332 5108 3384 5160
rect 3700 5108 3752 5160
rect 6276 5244 6328 5296
rect 7012 5244 7064 5296
rect 7932 5287 7984 5296
rect 7932 5253 7941 5287
rect 7941 5253 7975 5287
rect 7975 5253 7984 5287
rect 7932 5244 7984 5253
rect 2596 4972 2648 5024
rect 5172 4972 5224 5024
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 6644 5151 6696 5160
rect 6644 5117 6653 5151
rect 6653 5117 6687 5151
rect 6687 5117 6696 5151
rect 6644 5108 6696 5117
rect 9128 5176 9180 5228
rect 10784 5312 10836 5364
rect 15476 5312 15528 5364
rect 9864 5244 9916 5296
rect 10692 5244 10744 5296
rect 10232 5108 10284 5160
rect 10508 5176 10560 5228
rect 11244 5176 11296 5228
rect 12532 5244 12584 5296
rect 13176 5244 13228 5296
rect 13452 5244 13504 5296
rect 11980 5219 12032 5228
rect 11980 5185 11989 5219
rect 11989 5185 12023 5219
rect 12023 5185 12032 5219
rect 11980 5176 12032 5185
rect 12164 5176 12216 5228
rect 12348 5176 12400 5228
rect 12440 5176 12492 5228
rect 13360 5176 13412 5228
rect 15844 5176 15896 5228
rect 6828 5040 6880 5092
rect 9864 5040 9916 5092
rect 9956 5040 10008 5092
rect 10324 5040 10376 5092
rect 10600 5040 10652 5092
rect 10784 5108 10836 5160
rect 14004 5108 14056 5160
rect 11888 5040 11940 5092
rect 8668 4972 8720 5024
rect 8944 4972 8996 5024
rect 12348 5040 12400 5092
rect 12808 5040 12860 5092
rect 12256 4972 12308 5024
rect 12900 4972 12952 5024
rect 12992 4972 13044 5024
rect 14280 4972 14332 5024
rect 15200 5015 15252 5024
rect 15200 4981 15209 5015
rect 15209 4981 15243 5015
rect 15243 4981 15252 5015
rect 15200 4972 15252 4981
rect 15292 4972 15344 5024
rect 15476 4972 15528 5024
rect 2924 4870 2976 4922
rect 2988 4870 3040 4922
rect 3052 4870 3104 4922
rect 3116 4870 3168 4922
rect 3180 4870 3232 4922
rect 6872 4870 6924 4922
rect 6936 4870 6988 4922
rect 7000 4870 7052 4922
rect 7064 4870 7116 4922
rect 7128 4870 7180 4922
rect 10820 4870 10872 4922
rect 10884 4870 10936 4922
rect 10948 4870 11000 4922
rect 11012 4870 11064 4922
rect 11076 4870 11128 4922
rect 14768 4870 14820 4922
rect 14832 4870 14884 4922
rect 14896 4870 14948 4922
rect 14960 4870 15012 4922
rect 15024 4870 15076 4922
rect 1768 4768 1820 4820
rect 3148 4768 3200 4820
rect 3792 4768 3844 4820
rect 2596 4743 2648 4752
rect 2596 4709 2605 4743
rect 2605 4709 2639 4743
rect 2639 4709 2648 4743
rect 2596 4700 2648 4709
rect 4252 4768 4304 4820
rect 5080 4768 5132 4820
rect 7840 4768 7892 4820
rect 1492 4675 1544 4684
rect 1492 4641 1501 4675
rect 1501 4641 1535 4675
rect 1535 4641 1544 4675
rect 1492 4632 1544 4641
rect 1768 4564 1820 4616
rect 2228 4564 2280 4616
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 4068 4700 4120 4752
rect 3240 4632 3292 4684
rect 8300 4743 8352 4752
rect 8300 4709 8309 4743
rect 8309 4709 8343 4743
rect 8343 4709 8352 4743
rect 8944 4743 8996 4752
rect 8300 4700 8352 4709
rect 8944 4709 8953 4743
rect 8953 4709 8987 4743
rect 8987 4709 8996 4743
rect 8944 4700 8996 4709
rect 9128 4700 9180 4752
rect 9864 4768 9916 4820
rect 12072 4768 12124 4820
rect 12992 4811 13044 4820
rect 12992 4777 13001 4811
rect 13001 4777 13035 4811
rect 13035 4777 13044 4811
rect 12992 4768 13044 4777
rect 14280 4811 14332 4820
rect 14280 4777 14289 4811
rect 14289 4777 14323 4811
rect 14323 4777 14332 4811
rect 14280 4768 14332 4777
rect 3148 4607 3200 4616
rect 3148 4573 3157 4607
rect 3157 4573 3191 4607
rect 3191 4573 3200 4607
rect 3148 4564 3200 4573
rect 3332 4564 3384 4616
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 8024 4632 8076 4684
rect 8668 4632 8720 4684
rect 9496 4632 9548 4684
rect 10416 4700 10468 4752
rect 12348 4700 12400 4752
rect 12808 4700 12860 4752
rect 15936 4811 15988 4820
rect 15936 4777 15945 4811
rect 15945 4777 15979 4811
rect 15979 4777 15988 4811
rect 15936 4768 15988 4777
rect 14924 4700 14976 4752
rect 12532 4632 12584 4684
rect 9128 4607 9180 4616
rect 5816 4496 5868 4548
rect 6552 4496 6604 4548
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 10232 4564 10284 4616
rect 10784 4564 10836 4616
rect 10968 4564 11020 4616
rect 12808 4564 12860 4616
rect 13360 4564 13412 4616
rect 6736 4428 6788 4480
rect 8024 4428 8076 4480
rect 9772 4496 9824 4548
rect 8852 4428 8904 4480
rect 9128 4428 9180 4480
rect 11244 4428 11296 4480
rect 12256 4496 12308 4548
rect 12900 4496 12952 4548
rect 14648 4496 14700 4548
rect 14740 4496 14792 4548
rect 13452 4428 13504 4480
rect 14464 4471 14516 4480
rect 14464 4437 14473 4471
rect 14473 4437 14507 4471
rect 14507 4437 14516 4471
rect 14464 4428 14516 4437
rect 4898 4326 4950 4378
rect 4962 4326 5014 4378
rect 5026 4326 5078 4378
rect 5090 4326 5142 4378
rect 5154 4326 5206 4378
rect 8846 4326 8898 4378
rect 8910 4326 8962 4378
rect 8974 4326 9026 4378
rect 9038 4326 9090 4378
rect 9102 4326 9154 4378
rect 12794 4326 12846 4378
rect 12858 4326 12910 4378
rect 12922 4326 12974 4378
rect 12986 4326 13038 4378
rect 13050 4326 13102 4378
rect 2504 4224 2556 4276
rect 6460 4224 6512 4276
rect 9496 4224 9548 4276
rect 9772 4224 9824 4276
rect 10968 4224 11020 4276
rect 11060 4224 11112 4276
rect 12440 4224 12492 4276
rect 14464 4224 14516 4276
rect 14832 4224 14884 4276
rect 16764 4224 16816 4276
rect 1952 4156 2004 4208
rect 2412 4156 2464 4208
rect 2872 4199 2924 4208
rect 2872 4165 2906 4199
rect 2906 4165 2924 4199
rect 2872 4156 2924 4165
rect 2504 4088 2556 4140
rect 4436 4131 4488 4140
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 664 4020 716 4072
rect 2596 4063 2648 4072
rect 2228 3952 2280 4004
rect 2320 3884 2372 3936
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 6920 4088 6972 4140
rect 3792 3952 3844 4004
rect 5540 3952 5592 4004
rect 5724 3952 5776 4004
rect 6828 4020 6880 4072
rect 6368 3995 6420 4004
rect 6368 3961 6377 3995
rect 6377 3961 6411 3995
rect 6411 3961 6420 3995
rect 6368 3952 6420 3961
rect 7196 4088 7248 4140
rect 7380 4131 7432 4140
rect 7380 4097 7414 4131
rect 7414 4097 7432 4131
rect 7380 4088 7432 4097
rect 8668 4156 8720 4208
rect 8944 4156 8996 4208
rect 11520 4156 11572 4208
rect 11612 4156 11664 4208
rect 8852 4088 8904 4140
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 9680 4088 9732 4140
rect 11796 4156 11848 4208
rect 12164 4156 12216 4208
rect 12256 4156 12308 4208
rect 8484 4020 8536 4072
rect 8668 4020 8720 4072
rect 9496 4020 9548 4072
rect 9772 4020 9824 4072
rect 10600 4020 10652 4072
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 11152 4020 11204 4072
rect 12072 4088 12124 4140
rect 12348 4088 12400 4140
rect 13268 4156 13320 4208
rect 13728 4156 13780 4208
rect 14924 4156 14976 4208
rect 15936 4156 15988 4208
rect 13544 4088 13596 4140
rect 14096 4131 14148 4140
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 14096 4088 14148 4097
rect 14464 4088 14516 4140
rect 14832 4088 14884 4140
rect 16028 4131 16080 4140
rect 12164 4020 12216 4072
rect 13452 4020 13504 4072
rect 6092 3884 6144 3936
rect 8208 3952 8260 4004
rect 6644 3884 6696 3936
rect 8300 3884 8352 3936
rect 8484 3927 8536 3936
rect 8484 3893 8493 3927
rect 8493 3893 8527 3927
rect 8527 3893 8536 3927
rect 8484 3884 8536 3893
rect 8852 3884 8904 3936
rect 12256 3884 12308 3936
rect 14372 4020 14424 4072
rect 15108 4020 15160 4072
rect 16028 4097 16037 4131
rect 16037 4097 16071 4131
rect 16071 4097 16080 4131
rect 16028 4088 16080 4097
rect 16856 4020 16908 4072
rect 14740 3952 14792 4004
rect 14280 3884 14332 3936
rect 14556 3884 14608 3936
rect 15292 3884 15344 3936
rect 2924 3782 2976 3834
rect 2988 3782 3040 3834
rect 3052 3782 3104 3834
rect 3116 3782 3168 3834
rect 3180 3782 3232 3834
rect 6872 3782 6924 3834
rect 6936 3782 6988 3834
rect 7000 3782 7052 3834
rect 7064 3782 7116 3834
rect 7128 3782 7180 3834
rect 10820 3782 10872 3834
rect 10884 3782 10936 3834
rect 10948 3782 11000 3834
rect 11012 3782 11064 3834
rect 11076 3782 11128 3834
rect 14768 3782 14820 3834
rect 14832 3782 14884 3834
rect 14896 3782 14948 3834
rect 14960 3782 15012 3834
rect 15024 3782 15076 3834
rect 3516 3680 3568 3732
rect 6092 3680 6144 3732
rect 6184 3680 6236 3732
rect 6644 3680 6696 3732
rect 7104 3680 7156 3732
rect 10968 3723 11020 3732
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 2504 3544 2556 3596
rect 4160 3612 4212 3664
rect 4712 3612 4764 3664
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 3332 3476 3384 3528
rect 3516 3476 3568 3528
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 4252 3544 4304 3596
rect 4528 3544 4580 3596
rect 7196 3612 7248 3664
rect 6552 3544 6604 3596
rect 10968 3689 10977 3723
rect 10977 3689 11011 3723
rect 11011 3689 11020 3723
rect 10968 3680 11020 3689
rect 11888 3680 11940 3732
rect 12256 3680 12308 3732
rect 12348 3680 12400 3732
rect 14280 3723 14332 3732
rect 14280 3689 14289 3723
rect 14289 3689 14323 3723
rect 14323 3689 14332 3723
rect 14280 3680 14332 3689
rect 14556 3680 14608 3732
rect 16488 3680 16540 3732
rect 8024 3655 8076 3664
rect 8024 3621 8033 3655
rect 8033 3621 8067 3655
rect 8067 3621 8076 3655
rect 8024 3612 8076 3621
rect 9956 3612 10008 3664
rect 11704 3655 11756 3664
rect 11704 3621 11713 3655
rect 11713 3621 11747 3655
rect 11747 3621 11756 3655
rect 11704 3612 11756 3621
rect 12164 3612 12216 3664
rect 15752 3612 15804 3664
rect 8944 3587 8996 3596
rect 5448 3476 5500 3528
rect 6460 3476 6512 3528
rect 7288 3476 7340 3528
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 10232 3544 10284 3596
rect 940 3408 992 3460
rect 3700 3408 3752 3460
rect 6184 3408 6236 3460
rect 2872 3340 2924 3392
rect 7380 3408 7432 3460
rect 7748 3451 7800 3460
rect 7748 3417 7757 3451
rect 7757 3417 7791 3451
rect 7791 3417 7800 3451
rect 7748 3408 7800 3417
rect 8116 3476 8168 3528
rect 9496 3476 9548 3528
rect 11060 3544 11112 3596
rect 8208 3408 8260 3460
rect 7564 3340 7616 3392
rect 11244 3476 11296 3528
rect 11428 3476 11480 3528
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 12164 3476 12216 3528
rect 12256 3476 12308 3528
rect 12716 3519 12768 3528
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 12716 3476 12768 3485
rect 10784 3451 10836 3460
rect 10784 3417 10793 3451
rect 10793 3417 10827 3451
rect 10827 3417 10836 3451
rect 10784 3408 10836 3417
rect 10876 3408 10928 3460
rect 11152 3383 11204 3392
rect 11152 3349 11161 3383
rect 11161 3349 11195 3383
rect 11195 3349 11204 3383
rect 11520 3408 11572 3460
rect 11980 3408 12032 3460
rect 13176 3408 13228 3460
rect 13728 3408 13780 3460
rect 11152 3340 11204 3349
rect 13636 3340 13688 3392
rect 13912 3476 13964 3528
rect 16120 3476 16172 3528
rect 14464 3408 14516 3460
rect 16304 3340 16356 3392
rect 4898 3238 4950 3290
rect 4962 3238 5014 3290
rect 5026 3238 5078 3290
rect 5090 3238 5142 3290
rect 5154 3238 5206 3290
rect 8846 3238 8898 3290
rect 8910 3238 8962 3290
rect 8974 3238 9026 3290
rect 9038 3238 9090 3290
rect 9102 3238 9154 3290
rect 12794 3238 12846 3290
rect 12858 3238 12910 3290
rect 12922 3238 12974 3290
rect 12986 3238 13038 3290
rect 13050 3238 13102 3290
rect 2136 3136 2188 3188
rect 2504 3136 2556 3188
rect 4620 3136 4672 3188
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 5448 3068 5500 3120
rect 2872 3043 2924 3052
rect 2596 3000 2648 3009
rect 2872 3009 2906 3043
rect 2906 3009 2924 3043
rect 2872 3000 2924 3009
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 7012 3136 7064 3188
rect 7104 3136 7156 3188
rect 9772 3136 9824 3188
rect 9956 3136 10008 3188
rect 10508 3136 10560 3188
rect 10876 3136 10928 3188
rect 12072 3136 12124 3188
rect 12164 3136 12216 3188
rect 12532 3136 12584 3188
rect 13728 3136 13780 3188
rect 13820 3136 13872 3188
rect 15476 3136 15528 3188
rect 16488 3136 16540 3188
rect 6736 3111 6788 3120
rect 6736 3077 6745 3111
rect 6745 3077 6779 3111
rect 6779 3077 6788 3111
rect 6736 3068 6788 3077
rect 7472 3068 7524 3120
rect 8760 3068 8812 3120
rect 9036 3068 9088 3120
rect 9496 3068 9548 3120
rect 10048 3111 10100 3120
rect 10048 3077 10057 3111
rect 10057 3077 10091 3111
rect 10091 3077 10100 3111
rect 10048 3068 10100 3077
rect 11520 3111 11572 3120
rect 11520 3077 11529 3111
rect 11529 3077 11563 3111
rect 11563 3077 11572 3111
rect 11520 3068 11572 3077
rect 12440 3068 12492 3120
rect 13544 3068 13596 3120
rect 13912 3111 13964 3120
rect 13912 3077 13921 3111
rect 13921 3077 13955 3111
rect 13955 3077 13964 3111
rect 13912 3068 13964 3077
rect 14096 3111 14148 3120
rect 14096 3077 14105 3111
rect 14105 3077 14139 3111
rect 14139 3077 14148 3111
rect 14096 3068 14148 3077
rect 1492 2932 1544 2984
rect 2504 2932 2556 2984
rect 5448 2932 5500 2984
rect 5724 2932 5776 2984
rect 1952 2864 2004 2916
rect 2136 2864 2188 2916
rect 4160 2864 4212 2916
rect 5540 2864 5592 2916
rect 7564 2932 7616 2984
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 8668 2932 8720 2984
rect 9312 2932 9364 2984
rect 9772 3000 9824 3052
rect 12532 3000 12584 3052
rect 12716 3000 12768 3052
rect 13084 3000 13136 3052
rect 13268 3000 13320 3052
rect 13728 3000 13780 3052
rect 14372 3000 14424 3052
rect 11060 2932 11112 2984
rect 13544 2932 13596 2984
rect 14556 3000 14608 3052
rect 15384 3000 15436 3052
rect 15844 3000 15896 3052
rect 14740 2932 14792 2984
rect 8024 2864 8076 2916
rect 9680 2864 9732 2916
rect 12808 2864 12860 2916
rect 15108 2864 15160 2916
rect 4068 2796 4120 2848
rect 5172 2796 5224 2848
rect 8392 2796 8444 2848
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 10508 2796 10560 2848
rect 10784 2796 10836 2848
rect 11244 2796 11296 2848
rect 11888 2796 11940 2848
rect 12348 2796 12400 2848
rect 13084 2796 13136 2848
rect 13728 2796 13780 2848
rect 13820 2796 13872 2848
rect 14648 2839 14700 2848
rect 14648 2805 14657 2839
rect 14657 2805 14691 2839
rect 14691 2805 14700 2839
rect 14648 2796 14700 2805
rect 2924 2694 2976 2746
rect 2988 2694 3040 2746
rect 3052 2694 3104 2746
rect 3116 2694 3168 2746
rect 3180 2694 3232 2746
rect 6872 2694 6924 2746
rect 6936 2694 6988 2746
rect 7000 2694 7052 2746
rect 7064 2694 7116 2746
rect 7128 2694 7180 2746
rect 10820 2694 10872 2746
rect 10884 2694 10936 2746
rect 10948 2694 11000 2746
rect 11012 2694 11064 2746
rect 11076 2694 11128 2746
rect 14768 2694 14820 2746
rect 14832 2694 14884 2746
rect 14896 2694 14948 2746
rect 14960 2694 15012 2746
rect 15024 2694 15076 2746
rect 2780 2592 2832 2644
rect 3148 2592 3200 2644
rect 7840 2592 7892 2644
rect 8024 2635 8076 2644
rect 8024 2601 8033 2635
rect 8033 2601 8067 2635
rect 8067 2601 8076 2635
rect 8024 2592 8076 2601
rect 8208 2592 8260 2644
rect 10140 2592 10192 2644
rect 10692 2592 10744 2644
rect 11888 2592 11940 2644
rect 2136 2524 2188 2576
rect 4068 2524 4120 2576
rect 1768 2456 1820 2508
rect 2688 2456 2740 2508
rect 5908 2524 5960 2576
rect 8300 2524 8352 2576
rect 8852 2524 8904 2576
rect 11060 2524 11112 2576
rect 11980 2524 12032 2576
rect 12532 2524 12584 2576
rect 14188 2592 14240 2644
rect 15568 2592 15620 2644
rect 16212 2592 16264 2644
rect 14924 2524 14976 2576
rect 16488 2524 16540 2576
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 6184 2456 6236 2508
rect 5632 2388 5684 2440
rect 5724 2388 5776 2440
rect 6644 2388 6696 2440
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 7564 2388 7616 2440
rect 8668 2388 8720 2440
rect 9036 2388 9088 2440
rect 9220 2388 9272 2440
rect 9864 2388 9916 2440
rect 10600 2320 10652 2372
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 11612 2431 11664 2440
rect 11612 2397 11621 2431
rect 11621 2397 11655 2431
rect 11655 2397 11664 2431
rect 11612 2388 11664 2397
rect 12072 2456 12124 2508
rect 12164 2456 12216 2508
rect 12440 2456 12492 2508
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 12624 2456 12676 2508
rect 16580 2456 16632 2508
rect 11796 2388 11848 2397
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 12992 2388 13044 2440
rect 13084 2388 13136 2440
rect 13636 2388 13688 2440
rect 14188 2431 14240 2440
rect 14188 2397 14197 2431
rect 14197 2397 14231 2431
rect 14231 2397 14240 2431
rect 14188 2388 14240 2397
rect 14924 2388 14976 2440
rect 15200 2388 15252 2440
rect 15752 2388 15804 2440
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 3976 2252 4028 2304
rect 4436 2252 4488 2304
rect 4620 2252 4672 2304
rect 8852 2252 8904 2304
rect 9220 2252 9272 2304
rect 9496 2252 9548 2304
rect 10048 2252 10100 2304
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10232 2252 10284 2261
rect 10968 2252 11020 2304
rect 11060 2252 11112 2304
rect 12440 2252 12492 2304
rect 12808 2252 12860 2304
rect 12900 2252 12952 2304
rect 14832 2295 14884 2304
rect 14832 2261 14841 2295
rect 14841 2261 14875 2295
rect 14875 2261 14884 2295
rect 14832 2252 14884 2261
rect 4898 2150 4950 2202
rect 4962 2150 5014 2202
rect 5026 2150 5078 2202
rect 5090 2150 5142 2202
rect 5154 2150 5206 2202
rect 8846 2150 8898 2202
rect 8910 2150 8962 2202
rect 8974 2150 9026 2202
rect 9038 2150 9090 2202
rect 9102 2150 9154 2202
rect 12794 2150 12846 2202
rect 12858 2150 12910 2202
rect 12922 2150 12974 2202
rect 12986 2150 13038 2202
rect 13050 2150 13102 2202
rect 1032 1980 1084 2032
rect 3424 1980 3476 2032
rect 4160 2023 4212 2032
rect 4160 1989 4169 2023
rect 4169 1989 4203 2023
rect 4203 1989 4212 2023
rect 4160 1980 4212 1989
rect 4804 1980 4856 2032
rect 2228 1912 2280 1964
rect 4252 1955 4304 1964
rect 4252 1921 4261 1955
rect 4261 1921 4295 1955
rect 4295 1921 4304 1955
rect 4252 1912 4304 1921
rect 5172 1912 5224 1964
rect 5540 1955 5592 1964
rect 1952 1887 2004 1896
rect 1952 1853 1961 1887
rect 1961 1853 1995 1887
rect 1995 1853 2004 1887
rect 1952 1844 2004 1853
rect 2688 1887 2740 1896
rect 2688 1853 2697 1887
rect 2697 1853 2731 1887
rect 2731 1853 2740 1887
rect 2688 1844 2740 1853
rect 4068 1844 4120 1896
rect 5080 1844 5132 1896
rect 5540 1921 5549 1955
rect 5549 1921 5583 1955
rect 5583 1921 5592 1955
rect 5540 1912 5592 1921
rect 6000 2048 6052 2100
rect 9772 2048 9824 2100
rect 10048 2048 10100 2100
rect 6276 1980 6328 2032
rect 7012 1980 7064 2032
rect 3792 1776 3844 1828
rect 4252 1776 4304 1828
rect 6736 1912 6788 1964
rect 8576 1980 8628 2032
rect 9036 1980 9088 2032
rect 9680 1912 9732 1964
rect 9864 1955 9916 1964
rect 9864 1921 9873 1955
rect 9873 1921 9907 1955
rect 9907 1921 9916 1955
rect 9864 1912 9916 1921
rect 10232 2023 10284 2032
rect 10232 1989 10241 2023
rect 10241 1989 10275 2023
rect 10275 1989 10284 2023
rect 10232 1980 10284 1989
rect 2780 1708 2832 1760
rect 3332 1708 3384 1760
rect 7104 1776 7156 1828
rect 8300 1776 8352 1828
rect 8576 1776 8628 1828
rect 9772 1844 9824 1896
rect 11888 2048 11940 2100
rect 12072 2048 12124 2100
rect 10876 2023 10928 2032
rect 10876 1989 10885 2023
rect 10885 1989 10919 2023
rect 10919 1989 10928 2023
rect 10876 1980 10928 1989
rect 11336 1980 11388 2032
rect 12164 1980 12216 2032
rect 12808 1980 12860 2032
rect 13268 1980 13320 2032
rect 10784 1955 10836 1964
rect 10784 1921 10793 1955
rect 10793 1921 10827 1955
rect 10827 1921 10836 1955
rect 10784 1912 10836 1921
rect 10692 1844 10744 1896
rect 11152 1912 11204 1964
rect 11888 1955 11940 1964
rect 11336 1844 11388 1896
rect 11888 1921 11897 1955
rect 11897 1921 11931 1955
rect 11931 1921 11940 1955
rect 11888 1912 11940 1921
rect 12348 1955 12400 1964
rect 12348 1921 12357 1955
rect 12357 1921 12391 1955
rect 12391 1921 12400 1955
rect 12348 1912 12400 1921
rect 12440 1955 12492 1964
rect 12440 1921 12449 1955
rect 12449 1921 12483 1955
rect 12483 1921 12492 1955
rect 12440 1912 12492 1921
rect 12624 1912 12676 1964
rect 13728 2048 13780 2100
rect 15476 2048 15528 2100
rect 14004 2023 14056 2032
rect 14004 1989 14013 2023
rect 14013 1989 14047 2023
rect 14047 1989 14056 2023
rect 14004 1980 14056 1989
rect 14464 1980 14516 2032
rect 15016 1955 15068 1964
rect 15016 1921 15025 1955
rect 15025 1921 15059 1955
rect 15059 1921 15068 1955
rect 15016 1912 15068 1921
rect 9128 1708 9180 1760
rect 9312 1708 9364 1760
rect 10508 1776 10560 1828
rect 11796 1844 11848 1896
rect 13084 1844 13136 1896
rect 14096 1844 14148 1896
rect 12072 1776 12124 1828
rect 12164 1776 12216 1828
rect 13452 1776 13504 1828
rect 13728 1776 13780 1828
rect 10968 1708 11020 1760
rect 12992 1708 13044 1760
rect 13544 1708 13596 1760
rect 17316 1708 17368 1760
rect 2924 1606 2976 1658
rect 2988 1606 3040 1658
rect 3052 1606 3104 1658
rect 3116 1606 3168 1658
rect 3180 1606 3232 1658
rect 6872 1606 6924 1658
rect 6936 1606 6988 1658
rect 7000 1606 7052 1658
rect 7064 1606 7116 1658
rect 7128 1606 7180 1658
rect 10820 1606 10872 1658
rect 10884 1606 10936 1658
rect 10948 1606 11000 1658
rect 11012 1606 11064 1658
rect 11076 1606 11128 1658
rect 14768 1606 14820 1658
rect 14832 1606 14884 1658
rect 14896 1606 14948 1658
rect 14960 1606 15012 1658
rect 15024 1606 15076 1658
rect 1676 1504 1728 1556
rect 3240 1436 3292 1488
rect 4528 1436 4580 1488
rect 4712 1436 4764 1488
rect 5080 1504 5132 1556
rect 6460 1504 6512 1556
rect 6736 1504 6788 1556
rect 5448 1436 5500 1488
rect 6368 1436 6420 1488
rect 6644 1436 6696 1488
rect 8484 1504 8536 1556
rect 8944 1547 8996 1556
rect 8944 1513 8953 1547
rect 8953 1513 8987 1547
rect 8987 1513 8996 1547
rect 8944 1504 8996 1513
rect 9496 1504 9548 1556
rect 9956 1504 10008 1556
rect 10508 1504 10560 1556
rect 11520 1504 11572 1556
rect 11704 1547 11756 1556
rect 11704 1513 11713 1547
rect 11713 1513 11747 1547
rect 11747 1513 11756 1547
rect 11704 1504 11756 1513
rect 11796 1504 11848 1556
rect 12072 1504 12124 1556
rect 13268 1547 13320 1556
rect 9128 1436 9180 1488
rect 2044 1343 2096 1352
rect 2044 1309 2053 1343
rect 2053 1309 2087 1343
rect 2087 1309 2096 1343
rect 2044 1300 2096 1309
rect 572 1232 624 1284
rect 2320 1343 2372 1352
rect 2320 1309 2329 1343
rect 2329 1309 2363 1343
rect 2363 1309 2372 1343
rect 2320 1300 2372 1309
rect 756 1164 808 1216
rect 4252 1368 4304 1420
rect 4344 1368 4396 1420
rect 13268 1513 13277 1547
rect 13277 1513 13311 1547
rect 13311 1513 13320 1547
rect 13268 1504 13320 1513
rect 14188 1504 14240 1556
rect 14464 1547 14516 1556
rect 14464 1513 14473 1547
rect 14473 1513 14507 1547
rect 14507 1513 14516 1547
rect 14464 1504 14516 1513
rect 17408 1504 17460 1556
rect 13176 1436 13228 1488
rect 2964 1343 3016 1352
rect 2964 1309 2973 1343
rect 2973 1309 3007 1343
rect 3007 1309 3016 1343
rect 2964 1300 3016 1309
rect 3240 1343 3292 1352
rect 3240 1309 3249 1343
rect 3249 1309 3283 1343
rect 3283 1309 3292 1343
rect 3240 1300 3292 1309
rect 4068 1300 4120 1352
rect 3148 1207 3200 1216
rect 3148 1173 3157 1207
rect 3157 1173 3191 1207
rect 3191 1173 3200 1207
rect 3148 1164 3200 1173
rect 4620 1207 4672 1216
rect 4620 1173 4629 1207
rect 4629 1173 4663 1207
rect 4663 1173 4672 1207
rect 4620 1164 4672 1173
rect 5172 1300 5224 1352
rect 6644 1300 6696 1352
rect 6828 1343 6880 1352
rect 6828 1309 6837 1343
rect 6837 1309 6871 1343
rect 6871 1309 6880 1343
rect 6828 1300 6880 1309
rect 8392 1343 8444 1352
rect 8392 1309 8401 1343
rect 8401 1309 8435 1343
rect 8435 1309 8444 1343
rect 8392 1300 8444 1309
rect 8484 1300 8536 1352
rect 9036 1300 9088 1352
rect 6000 1232 6052 1284
rect 6552 1275 6604 1284
rect 6552 1241 6561 1275
rect 6561 1241 6595 1275
rect 6595 1241 6604 1275
rect 6552 1232 6604 1241
rect 8668 1232 8720 1284
rect 8944 1232 8996 1284
rect 9864 1275 9916 1284
rect 9864 1241 9873 1275
rect 9873 1241 9907 1275
rect 9907 1241 9916 1275
rect 9864 1232 9916 1241
rect 10508 1232 10560 1284
rect 7656 1164 7708 1216
rect 8116 1164 8168 1216
rect 10232 1207 10284 1216
rect 10232 1173 10241 1207
rect 10241 1173 10275 1207
rect 10275 1173 10284 1207
rect 10232 1164 10284 1173
rect 11244 1300 11296 1352
rect 11336 1300 11388 1352
rect 11428 1232 11480 1284
rect 11612 1300 11664 1352
rect 13636 1368 13688 1420
rect 12072 1232 12124 1284
rect 13268 1300 13320 1352
rect 13728 1300 13780 1352
rect 14280 1300 14332 1352
rect 15844 1343 15896 1352
rect 15844 1309 15853 1343
rect 15853 1309 15887 1343
rect 15887 1309 15896 1343
rect 15844 1300 15896 1309
rect 13084 1232 13136 1284
rect 11704 1207 11756 1216
rect 11704 1173 11729 1207
rect 11729 1173 11756 1207
rect 11704 1164 11756 1173
rect 13912 1232 13964 1284
rect 14096 1275 14148 1284
rect 14096 1241 14105 1275
rect 14105 1241 14139 1275
rect 14139 1241 14148 1275
rect 14096 1232 14148 1241
rect 13268 1164 13320 1216
rect 15660 1207 15712 1216
rect 15660 1173 15669 1207
rect 15669 1173 15703 1207
rect 15703 1173 15712 1207
rect 15660 1164 15712 1173
rect 4898 1062 4950 1114
rect 4962 1062 5014 1114
rect 5026 1062 5078 1114
rect 5090 1062 5142 1114
rect 5154 1062 5206 1114
rect 8846 1062 8898 1114
rect 8910 1062 8962 1114
rect 8974 1062 9026 1114
rect 9038 1062 9090 1114
rect 9102 1062 9154 1114
rect 12794 1062 12846 1114
rect 12858 1062 12910 1114
rect 12922 1062 12974 1114
rect 12986 1062 13038 1114
rect 13050 1062 13102 1114
rect 1216 960 1268 1012
rect 10416 960 10468 1012
rect 10508 960 10560 1012
rect 14464 960 14516 1012
rect 480 892 532 944
rect 8392 892 8444 944
rect 9864 892 9916 944
rect 14004 892 14056 944
rect 4620 824 4672 876
rect 16672 824 16724 876
rect 2780 756 2832 808
rect 8484 756 8536 808
rect 9588 756 9640 808
rect 15844 756 15896 808
rect 2320 688 2372 740
rect 5264 688 5316 740
rect 10324 688 10376 740
rect 9680 620 9732 672
rect 10232 620 10284 672
rect 16856 620 16908 672
rect 6644 552 6696 604
rect 10692 552 10744 604
rect 3976 484 4028 536
rect 11704 484 11756 536
rect 13360 484 13412 536
rect 4436 416 4488 468
rect 11336 416 11388 468
rect 6368 348 6420 400
rect 9404 348 9456 400
rect 16028 348 16080 400
rect 3240 280 3292 332
rect 13820 280 13872 332
rect 2228 212 2280 264
rect 9864 212 9916 264
rect 3148 144 3200 196
rect 11980 144 12032 196
rect 7748 8 7800 60
rect 15660 8 15712 60
<< metal2 >>
rect 1582 23216 1638 23225
rect 1582 23151 1638 23160
rect 1490 22536 1546 22545
rect 1490 22471 1492 22480
rect 1544 22471 1546 22480
rect 1492 22442 1544 22448
rect 1596 22234 1624 23151
rect 4898 22876 5206 22885
rect 4898 22874 4904 22876
rect 4960 22874 4984 22876
rect 5040 22874 5064 22876
rect 5120 22874 5144 22876
rect 5200 22874 5206 22876
rect 4960 22822 4962 22874
rect 5142 22822 5144 22874
rect 4898 22820 4904 22822
rect 4960 22820 4984 22822
rect 5040 22820 5064 22822
rect 5120 22820 5144 22822
rect 5200 22820 5206 22822
rect 4898 22811 5206 22820
rect 8846 22876 9154 22885
rect 8846 22874 8852 22876
rect 8908 22874 8932 22876
rect 8988 22874 9012 22876
rect 9068 22874 9092 22876
rect 9148 22874 9154 22876
rect 8908 22822 8910 22874
rect 9090 22822 9092 22874
rect 8846 22820 8852 22822
rect 8908 22820 8932 22822
rect 8988 22820 9012 22822
rect 9068 22820 9092 22822
rect 9148 22820 9154 22822
rect 8846 22811 9154 22820
rect 12794 22876 13102 22885
rect 12794 22874 12800 22876
rect 12856 22874 12880 22876
rect 12936 22874 12960 22876
rect 13016 22874 13040 22876
rect 13096 22874 13102 22876
rect 12856 22822 12858 22874
rect 13038 22822 13040 22874
rect 12794 22820 12800 22822
rect 12856 22820 12880 22822
rect 12936 22820 12960 22822
rect 13016 22820 13040 22822
rect 13096 22820 13102 22822
rect 12794 22811 13102 22820
rect 14188 22636 14240 22642
rect 14188 22578 14240 22584
rect 2924 22332 3232 22341
rect 2924 22330 2930 22332
rect 2986 22330 3010 22332
rect 3066 22330 3090 22332
rect 3146 22330 3170 22332
rect 3226 22330 3232 22332
rect 2986 22278 2988 22330
rect 3168 22278 3170 22330
rect 2924 22276 2930 22278
rect 2986 22276 3010 22278
rect 3066 22276 3090 22278
rect 3146 22276 3170 22278
rect 3226 22276 3232 22278
rect 2924 22267 3232 22276
rect 6872 22332 7180 22341
rect 6872 22330 6878 22332
rect 6934 22330 6958 22332
rect 7014 22330 7038 22332
rect 7094 22330 7118 22332
rect 7174 22330 7180 22332
rect 6934 22278 6936 22330
rect 7116 22278 7118 22330
rect 6872 22276 6878 22278
rect 6934 22276 6958 22278
rect 7014 22276 7038 22278
rect 7094 22276 7118 22278
rect 7174 22276 7180 22278
rect 6872 22267 7180 22276
rect 10820 22332 11128 22341
rect 10820 22330 10826 22332
rect 10882 22330 10906 22332
rect 10962 22330 10986 22332
rect 11042 22330 11066 22332
rect 11122 22330 11128 22332
rect 10882 22278 10884 22330
rect 11064 22278 11066 22330
rect 10820 22276 10826 22278
rect 10882 22276 10906 22278
rect 10962 22276 10986 22278
rect 11042 22276 11066 22278
rect 11122 22276 11128 22278
rect 10820 22267 11128 22276
rect 1584 22228 1636 22234
rect 1584 22170 1636 22176
rect 2780 22160 2832 22166
rect 2780 22102 2832 22108
rect 2410 21720 2466 21729
rect 388 21684 440 21690
rect 2410 21655 2466 21664
rect 388 21626 440 21632
rect 296 17876 348 17882
rect 296 17818 348 17824
rect 18 17776 74 17785
rect 18 17711 74 17720
rect 32 2553 60 17711
rect 308 12374 336 17818
rect 296 12368 348 12374
rect 296 12310 348 12316
rect 400 11558 428 21626
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1032 20460 1084 20466
rect 1032 20402 1084 20408
rect 478 19272 534 19281
rect 478 19207 534 19216
rect 492 12986 520 19207
rect 938 17640 994 17649
rect 938 17575 994 17584
rect 848 16788 900 16794
rect 848 16730 900 16736
rect 756 16448 808 16454
rect 756 16390 808 16396
rect 570 16280 626 16289
rect 570 16215 626 16224
rect 480 12980 532 12986
rect 480 12922 532 12928
rect 388 11552 440 11558
rect 388 11494 440 11500
rect 478 8256 534 8265
rect 478 8191 534 8200
rect 18 2544 74 2553
rect 18 2479 74 2488
rect 492 950 520 8191
rect 584 1290 612 16215
rect 662 15464 718 15473
rect 662 15399 718 15408
rect 676 4078 704 15399
rect 768 13938 796 16390
rect 756 13932 808 13938
rect 756 13874 808 13880
rect 754 13832 810 13841
rect 754 13767 810 13776
rect 664 4072 716 4078
rect 664 4014 716 4020
rect 572 1284 624 1290
rect 572 1226 624 1232
rect 768 1222 796 13767
rect 860 5302 888 16730
rect 952 12306 980 17575
rect 940 12300 992 12306
rect 940 12242 992 12248
rect 940 10464 992 10470
rect 940 10406 992 10412
rect 848 5296 900 5302
rect 848 5238 900 5244
rect 952 3466 980 10406
rect 1044 9722 1072 20402
rect 1308 18352 1360 18358
rect 1308 18294 1360 18300
rect 1124 17604 1176 17610
rect 1124 17546 1176 17552
rect 1136 14006 1164 17546
rect 1216 16108 1268 16114
rect 1216 16050 1268 16056
rect 1228 14278 1256 16050
rect 1216 14272 1268 14278
rect 1216 14214 1268 14220
rect 1216 14068 1268 14074
rect 1216 14010 1268 14016
rect 1124 14000 1176 14006
rect 1124 13942 1176 13948
rect 1124 12980 1176 12986
rect 1124 12922 1176 12928
rect 1032 9716 1084 9722
rect 1032 9658 1084 9664
rect 1032 8900 1084 8906
rect 1032 8842 1084 8848
rect 940 3460 992 3466
rect 940 3402 992 3408
rect 1044 2961 1072 8842
rect 1030 2952 1086 2961
rect 1030 2887 1086 2896
rect 1136 2774 1164 12922
rect 1044 2746 1164 2774
rect 1044 2038 1072 2746
rect 1032 2032 1084 2038
rect 1032 1974 1084 1980
rect 756 1216 808 1222
rect 756 1158 808 1164
rect 1228 1018 1256 14010
rect 1320 1465 1348 18294
rect 1412 15745 1440 21286
rect 2424 21146 2452 21655
rect 2412 21140 2464 21146
rect 2412 21082 2464 21088
rect 2792 20942 2820 22102
rect 8024 22092 8076 22098
rect 14200 22094 14228 22578
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 14768 22332 15076 22341
rect 14768 22330 14774 22332
rect 14830 22330 14854 22332
rect 14910 22330 14934 22332
rect 14990 22330 15014 22332
rect 15070 22330 15076 22332
rect 14830 22278 14832 22330
rect 15012 22278 15014 22330
rect 14768 22276 14774 22278
rect 14830 22276 14854 22278
rect 14910 22276 14934 22278
rect 14990 22276 15014 22278
rect 15070 22276 15076 22278
rect 14768 22267 15076 22276
rect 14200 22066 14412 22094
rect 8024 22034 8076 22040
rect 3884 22024 3936 22030
rect 3884 21966 3936 21972
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 2924 21244 3232 21253
rect 2924 21242 2930 21244
rect 2986 21242 3010 21244
rect 3066 21242 3090 21244
rect 3146 21242 3170 21244
rect 3226 21242 3232 21244
rect 2986 21190 2988 21242
rect 3168 21190 3170 21242
rect 2924 21188 2930 21190
rect 2986 21188 3010 21190
rect 3066 21188 3090 21190
rect 3146 21188 3170 21190
rect 3226 21188 3232 21190
rect 2924 21179 3232 21188
rect 1492 20936 1544 20942
rect 1492 20878 1544 20884
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 1504 19514 1532 20878
rect 1584 20800 1636 20806
rect 1584 20742 1636 20748
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1504 16454 1532 19314
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1596 16130 1624 20742
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1860 20256 1912 20262
rect 1860 20198 1912 20204
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1504 16102 1624 16130
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1400 15632 1452 15638
rect 1400 15574 1452 15580
rect 1412 15366 1440 15574
rect 1400 15360 1452 15366
rect 1400 15302 1452 15308
rect 1412 14346 1440 15302
rect 1400 14340 1452 14346
rect 1400 14282 1452 14288
rect 1504 14249 1532 16102
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1596 15026 1624 15982
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1584 14884 1636 14890
rect 1584 14826 1636 14832
rect 1596 14482 1624 14826
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1584 14340 1636 14346
rect 1584 14282 1636 14288
rect 1490 14240 1546 14249
rect 1490 14175 1546 14184
rect 1400 14000 1452 14006
rect 1400 13942 1452 13948
rect 1412 10198 1440 13942
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1504 13326 1532 13670
rect 1596 13433 1624 14282
rect 1582 13424 1638 13433
rect 1582 13359 1638 13368
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1400 10192 1452 10198
rect 1400 10134 1452 10140
rect 1504 10130 1532 13262
rect 1582 13016 1638 13025
rect 1582 12951 1638 12960
rect 1596 11762 1624 12951
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 10606 1624 10950
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1596 10010 1624 10542
rect 1412 9982 1624 10010
rect 1412 5234 1440 9982
rect 1584 9716 1636 9722
rect 1688 9704 1716 19314
rect 1780 18290 1808 20198
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 16522 1808 18226
rect 1768 16516 1820 16522
rect 1768 16458 1820 16464
rect 1780 14958 1808 16458
rect 1872 16130 1900 20198
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1964 17678 1992 18362
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 1964 17202 1992 17614
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1964 16425 1992 17138
rect 1950 16416 2006 16425
rect 1950 16351 2006 16360
rect 1872 16102 1992 16130
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1872 15162 1900 15982
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1780 14006 1808 14758
rect 1872 14618 1900 14962
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1768 14000 1820 14006
rect 1768 13942 1820 13948
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1780 10810 1808 13806
rect 1872 13530 1900 14214
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1858 13424 1914 13433
rect 1858 13359 1860 13368
rect 1912 13359 1914 13368
rect 1860 13330 1912 13336
rect 1872 11082 1900 13330
rect 1964 12753 1992 16102
rect 2056 13258 2084 19246
rect 2136 17264 2188 17270
rect 2136 17206 2188 17212
rect 2148 15706 2176 17206
rect 2240 16250 2268 20878
rect 2688 20868 2740 20874
rect 2688 20810 2740 20816
rect 2412 20324 2464 20330
rect 2412 20266 2464 20272
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2332 19378 2360 20198
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2240 16017 2268 16050
rect 2226 16008 2282 16017
rect 2226 15943 2282 15952
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2332 15552 2360 18702
rect 2424 16561 2452 20266
rect 2700 19666 2728 20810
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2792 20233 2820 20538
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3160 20369 3188 20402
rect 3332 20392 3384 20398
rect 3146 20360 3202 20369
rect 3332 20334 3384 20340
rect 3146 20295 3202 20304
rect 2778 20224 2834 20233
rect 2778 20159 2834 20168
rect 2924 20156 3232 20165
rect 2924 20154 2930 20156
rect 2986 20154 3010 20156
rect 3066 20154 3090 20156
rect 3146 20154 3170 20156
rect 3226 20154 3232 20156
rect 2986 20102 2988 20154
rect 3168 20102 3170 20154
rect 2924 20100 2930 20102
rect 2986 20100 3010 20102
rect 3066 20100 3090 20102
rect 3146 20100 3170 20102
rect 3226 20100 3232 20102
rect 2924 20091 3232 20100
rect 3146 19952 3202 19961
rect 3202 19910 3280 19938
rect 3146 19887 3202 19896
rect 2870 19816 2926 19825
rect 2870 19751 2872 19760
rect 2924 19751 2926 19760
rect 2872 19722 2924 19728
rect 2700 19638 2912 19666
rect 2596 19440 2648 19446
rect 2594 19408 2596 19417
rect 2688 19440 2740 19446
rect 2648 19408 2650 19417
rect 2688 19382 2740 19388
rect 2594 19343 2650 19352
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2608 18873 2636 19246
rect 2594 18864 2650 18873
rect 2594 18799 2650 18808
rect 2608 18630 2636 18799
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2700 18272 2728 19382
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2884 19334 2912 19638
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 2792 18902 2820 19314
rect 2884 19306 3004 19334
rect 2976 19156 3004 19306
rect 3160 19242 3188 19450
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 2853 19128 3004 19156
rect 3252 19156 3280 19910
rect 3344 19854 3372 20334
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3330 19680 3386 19689
rect 3330 19615 3386 19624
rect 3344 19281 3372 19615
rect 3330 19272 3386 19281
rect 3330 19207 3386 19216
rect 3252 19128 3372 19156
rect 2853 18952 2881 19128
rect 2924 19068 3232 19077
rect 2924 19066 2930 19068
rect 2986 19066 3010 19068
rect 3066 19066 3090 19068
rect 3146 19066 3170 19068
rect 3226 19066 3232 19068
rect 2986 19014 2988 19066
rect 3168 19014 3170 19066
rect 2924 19012 2930 19014
rect 2986 19012 3010 19014
rect 3066 19012 3090 19014
rect 3146 19012 3170 19014
rect 3226 19012 3232 19014
rect 2924 19003 3232 19012
rect 3344 18952 3372 19128
rect 2853 18924 2912 18952
rect 2780 18896 2832 18902
rect 2780 18838 2832 18844
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2516 18244 2728 18272
rect 2410 16552 2466 16561
rect 2410 16487 2466 16496
rect 2410 16416 2466 16425
rect 2410 16351 2466 16360
rect 2424 16250 2452 16351
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2516 16182 2544 18244
rect 2686 18184 2742 18193
rect 2686 18119 2742 18128
rect 2596 17604 2648 17610
rect 2596 17546 2648 17552
rect 2608 16590 2636 17546
rect 2596 16584 2648 16590
rect 2700 16561 2728 18119
rect 2596 16526 2648 16532
rect 2686 16552 2742 16561
rect 2504 16176 2556 16182
rect 2504 16118 2556 16124
rect 2608 16046 2636 16526
rect 2686 16487 2742 16496
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2608 15638 2636 15982
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2148 15524 2360 15552
rect 2504 15564 2556 15570
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2148 12986 2176 15524
rect 2504 15506 2556 15512
rect 2320 15428 2372 15434
rect 2320 15370 2372 15376
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2240 14006 2268 15098
rect 2332 15026 2360 15370
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2240 13394 2268 13670
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2332 13002 2360 14962
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2424 13938 2452 14214
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2412 13796 2464 13802
rect 2412 13738 2464 13744
rect 2424 13297 2452 13738
rect 2410 13288 2466 13297
rect 2410 13223 2466 13232
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2240 12974 2360 13002
rect 2240 12889 2268 12974
rect 2320 12912 2372 12918
rect 2226 12880 2282 12889
rect 2044 12844 2096 12850
rect 2320 12854 2372 12860
rect 2226 12815 2282 12824
rect 2044 12786 2096 12792
rect 1950 12744 2006 12753
rect 1950 12679 2006 12688
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1768 10804 1820 10810
rect 1820 10764 1900 10792
rect 1768 10746 1820 10752
rect 1766 10704 1822 10713
rect 1766 10639 1768 10648
rect 1820 10639 1822 10648
rect 1768 10610 1820 10616
rect 1688 9676 1808 9704
rect 1584 9658 1636 9664
rect 1596 9602 1624 9658
rect 1596 9574 1716 9602
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 6866 1532 7346
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1504 6322 1532 6802
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1504 5778 1532 6054
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1504 3233 1532 4626
rect 1490 3224 1546 3233
rect 1490 3159 1546 3168
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1306 1456 1362 1465
rect 1306 1391 1362 1400
rect 1504 1329 1532 2926
rect 1596 2774 1624 8366
rect 1688 4706 1716 9574
rect 1780 6866 1808 9676
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1872 5234 1900 10764
rect 1964 8090 1992 12582
rect 2056 12442 2084 12786
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 2148 12306 2176 12582
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2240 11914 2268 12718
rect 2332 12356 2360 12854
rect 2516 12714 2544 15506
rect 2700 15484 2728 16186
rect 2608 15456 2728 15484
rect 2608 14958 2636 15456
rect 2688 15088 2740 15094
rect 2688 15030 2740 15036
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2594 14648 2650 14657
rect 2594 14583 2650 14592
rect 2608 13938 2636 14583
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2700 13818 2728 15030
rect 2608 13790 2728 13818
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2332 12328 2544 12356
rect 2608 12345 2636 13790
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2410 12200 2466 12209
rect 2332 12073 2360 12174
rect 2410 12135 2466 12144
rect 2318 12064 2374 12073
rect 2318 11999 2374 12008
rect 2240 11886 2360 11914
rect 2226 11792 2282 11801
rect 2136 11756 2188 11762
rect 2226 11727 2282 11736
rect 2136 11698 2188 11704
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 2056 8294 2084 11494
rect 2148 10810 2176 11698
rect 2240 11694 2268 11727
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2240 10577 2268 11630
rect 2332 11558 2360 11886
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2226 10568 2282 10577
rect 2226 10503 2282 10512
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2136 9512 2188 9518
rect 2134 9480 2136 9489
rect 2188 9480 2190 9489
rect 2134 9415 2190 9424
rect 2332 9058 2360 9590
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2240 9030 2360 9058
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1964 7546 1992 8026
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1780 4826 1808 5102
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1688 4678 1900 4706
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1596 2746 1716 2774
rect 1688 1562 1716 2746
rect 1780 2514 1808 4558
rect 1872 2938 1900 4678
rect 1964 4214 1992 5306
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1964 3058 1992 3538
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1872 2922 1992 2938
rect 1872 2916 2004 2922
rect 1872 2910 1952 2916
rect 1952 2858 2004 2864
rect 1768 2508 1820 2514
rect 1768 2450 1820 2456
rect 1952 1896 2004 1902
rect 1952 1838 2004 1844
rect 1676 1556 1728 1562
rect 1676 1498 1728 1504
rect 1490 1320 1546 1329
rect 1490 1255 1546 1264
rect 1216 1012 1268 1018
rect 1216 954 1268 960
rect 480 944 532 950
rect 480 886 532 892
rect 1964 649 1992 1838
rect 2056 1358 2084 5510
rect 2148 3194 2176 8978
rect 2240 7002 2268 9030
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2332 8090 2360 8230
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2240 4622 2268 6938
rect 2318 6216 2374 6225
rect 2318 6151 2374 6160
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2332 4026 2360 6151
rect 2424 4622 2452 12135
rect 2516 7834 2544 12328
rect 2594 12336 2650 12345
rect 2594 12271 2650 12280
rect 2608 12238 2636 12271
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2700 12102 2728 12786
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2594 11928 2650 11937
rect 2792 11898 2820 18634
rect 2884 18290 2912 18924
rect 3252 18924 3372 18952
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 3068 18601 3096 18770
rect 3054 18592 3110 18601
rect 3054 18527 3110 18536
rect 3252 18426 3280 18924
rect 3240 18420 3292 18426
rect 3240 18362 3292 18368
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 3436 18170 3464 21286
rect 3620 20874 3648 21286
rect 3608 20868 3660 20874
rect 3608 20810 3660 20816
rect 3700 20800 3752 20806
rect 3700 20742 3752 20748
rect 3792 20800 3844 20806
rect 3792 20742 3844 20748
rect 3516 20324 3568 20330
rect 3516 20266 3568 20272
rect 3528 19990 3556 20266
rect 3606 20224 3662 20233
rect 3606 20159 3662 20168
rect 3516 19984 3568 19990
rect 3516 19926 3568 19932
rect 3528 19786 3556 19926
rect 3620 19922 3648 20159
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3516 19780 3568 19786
rect 3516 19722 3568 19728
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3516 19440 3568 19446
rect 3516 19382 3568 19388
rect 3344 18142 3464 18170
rect 2924 17980 3232 17989
rect 2924 17978 2930 17980
rect 2986 17978 3010 17980
rect 3066 17978 3090 17980
rect 3146 17978 3170 17980
rect 3226 17978 3232 17980
rect 2986 17926 2988 17978
rect 3168 17926 3170 17978
rect 2924 17924 2930 17926
rect 2986 17924 3010 17926
rect 3066 17924 3090 17926
rect 3146 17924 3170 17926
rect 3226 17924 3232 17926
rect 2924 17915 3232 17924
rect 3344 17241 3372 18142
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3330 17232 3386 17241
rect 2964 17196 3016 17202
rect 3330 17167 3386 17176
rect 2964 17138 3016 17144
rect 2976 16980 3004 17138
rect 2853 16952 3004 16980
rect 2853 16776 2881 16952
rect 2924 16892 3232 16901
rect 2924 16890 2930 16892
rect 2986 16890 3010 16892
rect 3066 16890 3090 16892
rect 3146 16890 3170 16892
rect 3226 16890 3232 16892
rect 2986 16838 2988 16890
rect 3168 16838 3170 16890
rect 2924 16836 2930 16838
rect 2986 16836 3010 16838
rect 3066 16836 3090 16838
rect 3146 16836 3170 16838
rect 3226 16836 3232 16838
rect 2924 16827 3232 16836
rect 2853 16748 2912 16776
rect 2884 16182 2912 16748
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2884 15892 2912 16118
rect 2853 15864 2912 15892
rect 2853 15688 2881 15864
rect 2924 15804 3232 15813
rect 2924 15802 2930 15804
rect 2986 15802 3010 15804
rect 3066 15802 3090 15804
rect 3146 15802 3170 15804
rect 3226 15802 3232 15804
rect 2986 15750 2988 15802
rect 3168 15750 3170 15802
rect 2924 15748 2930 15750
rect 2986 15748 3010 15750
rect 3066 15748 3090 15750
rect 3146 15748 3170 15750
rect 3226 15748 3232 15750
rect 2924 15739 3232 15748
rect 2853 15660 3004 15688
rect 2976 15094 3004 15660
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 2872 15020 2924 15026
rect 2853 14968 2872 15008
rect 2853 14962 2924 14968
rect 2853 14600 2881 14962
rect 2924 14716 3232 14725
rect 2924 14714 2930 14716
rect 2986 14714 3010 14716
rect 3066 14714 3090 14716
rect 3146 14714 3170 14716
rect 3226 14714 3232 14716
rect 2986 14662 2988 14714
rect 3168 14662 3170 14714
rect 2924 14660 2930 14662
rect 2986 14660 3010 14662
rect 3066 14660 3090 14662
rect 3146 14660 3170 14662
rect 3226 14660 3232 14662
rect 2924 14651 3232 14660
rect 2853 14572 2912 14600
rect 2884 13734 2912 14572
rect 2964 13864 3016 13870
rect 2962 13832 2964 13841
rect 3016 13832 3018 13841
rect 2962 13767 3018 13776
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2924 13628 3232 13637
rect 2924 13626 2930 13628
rect 2986 13626 3010 13628
rect 3066 13626 3090 13628
rect 3146 13626 3170 13628
rect 3226 13626 3232 13628
rect 2986 13574 2988 13626
rect 3168 13574 3170 13626
rect 2924 13572 2930 13574
rect 2986 13572 3010 13574
rect 3066 13572 3090 13574
rect 3146 13572 3170 13574
rect 3226 13572 3232 13574
rect 2924 13563 3232 13572
rect 2872 13456 2924 13462
rect 2870 13424 2872 13433
rect 2924 13424 2926 13433
rect 2870 13359 2926 13368
rect 3146 13424 3202 13433
rect 3146 13359 3202 13368
rect 3240 13388 3292 13394
rect 3056 13320 3108 13326
rect 2976 13280 3056 13308
rect 2976 12764 3004 13280
rect 3056 13262 3108 13268
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 3068 12986 3096 13126
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3056 12776 3108 12782
rect 2976 12736 3056 12764
rect 3056 12718 3108 12724
rect 3160 12764 3188 13359
rect 3240 13330 3292 13336
rect 3252 13258 3280 13330
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3240 12776 3292 12782
rect 3160 12736 3240 12764
rect 3160 12628 3188 12736
rect 3240 12718 3292 12724
rect 2853 12600 3188 12628
rect 2853 12434 2881 12600
rect 2924 12540 3232 12549
rect 2924 12538 2930 12540
rect 2986 12538 3010 12540
rect 3066 12538 3090 12540
rect 3146 12538 3170 12540
rect 3226 12538 3232 12540
rect 2986 12486 2988 12538
rect 3168 12486 3170 12538
rect 2924 12484 2930 12486
rect 2986 12484 3010 12486
rect 3066 12484 3090 12486
rect 3146 12484 3170 12486
rect 3226 12484 3232 12486
rect 2924 12475 3232 12484
rect 3344 12434 3372 16390
rect 2853 12406 2912 12434
rect 2594 11863 2650 11872
rect 2780 11892 2832 11898
rect 2608 11014 2636 11863
rect 2780 11834 2832 11840
rect 2884 11608 2912 12406
rect 3252 12406 3372 12434
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2700 11580 2912 11608
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2594 10840 2650 10849
rect 2594 10775 2650 10784
rect 2608 7936 2636 10775
rect 2700 10606 2728 11580
rect 2976 11540 3004 11834
rect 3068 11626 3096 12310
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3160 11937 3188 12242
rect 3146 11928 3202 11937
rect 3146 11863 3202 11872
rect 3252 11762 3280 12406
rect 3436 12374 3464 18022
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3424 12232 3476 12238
rect 3422 12200 3424 12209
rect 3476 12200 3478 12209
rect 3422 12135 3478 12144
rect 3422 12064 3478 12073
rect 3422 11999 3478 12008
rect 3436 11898 3464 11999
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3528 11778 3556 19382
rect 3620 12617 3648 19654
rect 3712 18737 3740 20742
rect 3804 20097 3832 20742
rect 3790 20088 3846 20097
rect 3790 20023 3846 20032
rect 3792 19984 3844 19990
rect 3792 19926 3844 19932
rect 3698 18728 3754 18737
rect 3804 18698 3832 19926
rect 3896 18902 3924 21966
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 4898 21788 5206 21797
rect 4898 21786 4904 21788
rect 4960 21786 4984 21788
rect 5040 21786 5064 21788
rect 5120 21786 5144 21788
rect 5200 21786 5206 21788
rect 4960 21734 4962 21786
rect 5142 21734 5144 21786
rect 4898 21732 4904 21734
rect 4960 21732 4984 21734
rect 5040 21732 5064 21734
rect 5120 21732 5144 21734
rect 5200 21732 5206 21734
rect 4898 21723 5206 21732
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3988 20058 4016 20878
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 3974 19952 4030 19961
rect 3974 19887 4030 19896
rect 3988 19718 4016 19887
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3884 18896 3936 18902
rect 3884 18838 3936 18844
rect 3976 18896 4028 18902
rect 4080 18873 4108 21422
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4172 20466 4200 20742
rect 4898 20700 5206 20709
rect 4898 20698 4904 20700
rect 4960 20698 4984 20700
rect 5040 20698 5064 20700
rect 5120 20698 5144 20700
rect 5200 20698 5206 20700
rect 4960 20646 4962 20698
rect 5142 20646 5144 20698
rect 4898 20644 4904 20646
rect 4960 20644 4984 20646
rect 5040 20644 5064 20646
rect 5120 20644 5144 20646
rect 5200 20644 5206 20646
rect 4898 20635 5206 20644
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 4172 19922 4200 20266
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 3976 18838 4028 18844
rect 4066 18864 4122 18873
rect 3698 18663 3754 18672
rect 3792 18692 3844 18698
rect 3792 18634 3844 18640
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3790 18456 3846 18465
rect 3790 18391 3846 18400
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3712 17542 3740 18226
rect 3804 18222 3832 18391
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3804 17202 3832 18158
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3712 13462 3740 15846
rect 3804 15638 3832 17138
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3804 13172 3832 15438
rect 3896 13569 3924 18566
rect 3988 16182 4016 18838
rect 4066 18799 4122 18808
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 4080 18193 4108 18634
rect 4066 18184 4122 18193
rect 4066 18119 4122 18128
rect 4068 18080 4120 18086
rect 4066 18048 4068 18057
rect 4120 18048 4122 18057
rect 4066 17983 4122 17992
rect 4172 17678 4200 19450
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3974 16008 4030 16017
rect 3974 15943 4030 15952
rect 3988 15706 4016 15943
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3988 14056 4016 15302
rect 4080 14249 4108 16458
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 4172 14958 4200 15574
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4066 14240 4122 14249
rect 4066 14175 4122 14184
rect 3988 14028 4108 14056
rect 3974 13968 4030 13977
rect 3974 13903 3976 13912
rect 4028 13903 4030 13912
rect 3976 13874 4028 13880
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3882 13560 3938 13569
rect 3882 13495 3938 13504
rect 3712 13144 3832 13172
rect 3882 13152 3938 13161
rect 3712 12822 3740 13144
rect 3882 13087 3938 13096
rect 3712 12794 3832 12822
rect 3698 12744 3754 12753
rect 3698 12679 3754 12688
rect 3606 12608 3662 12617
rect 3606 12543 3662 12552
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3436 11750 3556 11778
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 2792 11512 3004 11540
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2700 8673 2728 10542
rect 2792 9994 2820 11512
rect 2924 11452 3232 11461
rect 2924 11450 2930 11452
rect 2986 11450 3010 11452
rect 3066 11450 3090 11452
rect 3146 11450 3170 11452
rect 3226 11450 3232 11452
rect 2986 11398 2988 11450
rect 3168 11398 3170 11450
rect 2924 11396 2930 11398
rect 2986 11396 3010 11398
rect 3066 11396 3090 11398
rect 3146 11396 3170 11398
rect 3226 11396 3232 11398
rect 2924 11387 3232 11396
rect 2962 11248 3018 11257
rect 2962 11183 2964 11192
rect 3016 11183 3018 11192
rect 3436 11200 3464 11750
rect 3516 11620 3568 11626
rect 3620 11608 3648 12310
rect 3568 11580 3648 11608
rect 3516 11562 3568 11568
rect 3606 11384 3662 11393
rect 3606 11319 3662 11328
rect 3436 11172 3556 11200
rect 2964 11154 3016 11160
rect 2870 11112 2926 11121
rect 2870 11047 2926 11056
rect 3424 11076 3476 11082
rect 2884 10674 2912 11047
rect 3424 11018 3476 11024
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2924 10364 3232 10373
rect 2924 10362 2930 10364
rect 2986 10362 3010 10364
rect 3066 10362 3090 10364
rect 3146 10362 3170 10364
rect 3226 10362 3232 10364
rect 2986 10310 2988 10362
rect 3168 10310 3170 10362
rect 2924 10308 2930 10310
rect 2986 10308 3010 10310
rect 3066 10308 3090 10310
rect 3146 10308 3170 10310
rect 3226 10308 3232 10310
rect 2924 10299 3232 10308
rect 3146 10160 3202 10169
rect 3344 10112 3372 10950
rect 3146 10095 3148 10104
rect 3200 10095 3202 10104
rect 3148 10066 3200 10072
rect 3252 10084 3372 10112
rect 3146 10024 3202 10033
rect 2780 9988 2832 9994
rect 3146 9959 3202 9968
rect 2780 9930 2832 9936
rect 3160 9518 3188 9959
rect 3252 9586 3280 10084
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2686 8664 2742 8673
rect 2686 8599 2742 8608
rect 2608 7908 2728 7936
rect 2516 7806 2636 7834
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 4729 2544 7686
rect 2608 5370 2636 7806
rect 2700 7342 2728 7908
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2700 6905 2728 7278
rect 2686 6896 2742 6905
rect 2686 6831 2742 6840
rect 2792 6610 2820 9386
rect 2924 9276 3232 9285
rect 2924 9274 2930 9276
rect 2986 9274 3010 9276
rect 3066 9274 3090 9276
rect 3146 9274 3170 9276
rect 3226 9274 3232 9276
rect 2986 9222 2988 9274
rect 3168 9222 3170 9274
rect 2924 9220 2930 9222
rect 2986 9220 3010 9222
rect 3066 9220 3090 9222
rect 3146 9220 3170 9222
rect 3226 9220 3232 9222
rect 2924 9211 3232 9220
rect 2924 8188 3232 8197
rect 2924 8186 2930 8188
rect 2986 8186 3010 8188
rect 3066 8186 3090 8188
rect 3146 8186 3170 8188
rect 3226 8186 3232 8188
rect 2986 8134 2988 8186
rect 3168 8134 3170 8186
rect 2924 8132 2930 8134
rect 2986 8132 3010 8134
rect 3066 8132 3090 8134
rect 3146 8132 3170 8134
rect 3226 8132 3232 8134
rect 2924 8123 3232 8132
rect 3344 7750 3372 9930
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 2924 7100 3232 7109
rect 2924 7098 2930 7100
rect 2986 7098 3010 7100
rect 3066 7098 3090 7100
rect 3146 7098 3170 7100
rect 3226 7098 3232 7100
rect 2986 7046 2988 7098
rect 3168 7046 3170 7098
rect 2924 7044 2930 7046
rect 2986 7044 3010 7046
rect 3066 7044 3090 7046
rect 3146 7044 3170 7046
rect 3226 7044 3232 7046
rect 2924 7035 3232 7044
rect 2700 6582 2820 6610
rect 2700 5817 2728 6582
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2686 5808 2742 5817
rect 2686 5743 2742 5752
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2608 4758 2636 4966
rect 2596 4752 2648 4758
rect 2502 4720 2558 4729
rect 2596 4694 2648 4700
rect 2502 4655 2558 4664
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2516 4282 2544 4655
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2240 4010 2360 4026
rect 2228 4004 2360 4010
rect 2280 3998 2360 4004
rect 2228 3946 2280 3952
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2136 2916 2188 2922
rect 2136 2858 2188 2864
rect 2148 2582 2176 2858
rect 2136 2576 2188 2582
rect 2136 2518 2188 2524
rect 2228 1964 2280 1970
rect 2228 1906 2280 1912
rect 2044 1352 2096 1358
rect 2044 1294 2096 1300
rect 1950 640 2006 649
rect 1950 575 2006 584
rect 2240 270 2268 1906
rect 2332 1358 2360 3878
rect 2424 2774 2452 4150
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 3602 2544 4082
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2516 2990 2544 3130
rect 2608 3058 2636 4014
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2424 2746 2544 2774
rect 2516 2417 2544 2746
rect 2700 2514 2728 5743
rect 2792 5574 2820 6394
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 2924 6012 3232 6021
rect 2924 6010 2930 6012
rect 2986 6010 3010 6012
rect 3066 6010 3090 6012
rect 3146 6010 3170 6012
rect 3226 6010 3232 6012
rect 2986 5958 2988 6010
rect 3168 5958 3170 6010
rect 2924 5956 2930 5958
rect 2986 5956 3010 5958
rect 3066 5956 3090 5958
rect 3146 5956 3170 5958
rect 3226 5956 3232 5958
rect 2924 5947 3232 5956
rect 3344 5846 3372 6054
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 2792 4570 2820 5199
rect 3344 5166 3372 5646
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3330 4992 3386 5001
rect 2924 4924 3232 4933
rect 3330 4927 3386 4936
rect 2924 4922 2930 4924
rect 2986 4922 3010 4924
rect 3066 4922 3090 4924
rect 3146 4922 3170 4924
rect 3226 4922 3232 4924
rect 2986 4870 2988 4922
rect 3168 4870 3170 4922
rect 2924 4868 2930 4870
rect 2986 4868 3010 4870
rect 3066 4868 3090 4870
rect 3146 4868 3170 4870
rect 3226 4868 3232 4870
rect 2924 4859 3232 4868
rect 3148 4820 3200 4826
rect 3344 4808 3372 4927
rect 3148 4762 3200 4768
rect 3252 4780 3372 4808
rect 3160 4622 3188 4762
rect 3252 4690 3280 4780
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3148 4616 3200 4622
rect 2792 4542 3004 4570
rect 3148 4558 3200 4564
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 2870 4312 2926 4321
rect 2870 4247 2926 4256
rect 2884 4214 2912 4247
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2976 3924 3004 4542
rect 2792 3896 3004 3924
rect 2792 2650 2820 3896
rect 2924 3836 3232 3845
rect 2924 3834 2930 3836
rect 2986 3834 3010 3836
rect 3066 3834 3090 3836
rect 3146 3834 3170 3836
rect 3226 3834 3232 3836
rect 2986 3782 2988 3834
rect 3168 3782 3170 3834
rect 2924 3780 2930 3782
rect 2986 3780 3010 3782
rect 3066 3780 3090 3782
rect 3146 3780 3170 3782
rect 3226 3780 3232 3782
rect 2924 3771 3232 3780
rect 3344 3534 3372 4558
rect 3148 3528 3200 3534
rect 3146 3496 3148 3505
rect 3332 3528 3384 3534
rect 3200 3496 3202 3505
rect 3332 3470 3384 3476
rect 3146 3431 3202 3440
rect 2872 3392 2924 3398
rect 3436 3380 3464 11018
rect 3528 10441 3556 11172
rect 3514 10432 3570 10441
rect 3514 10367 3570 10376
rect 3620 8634 3648 11319
rect 3712 10674 3740 12679
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3606 8528 3662 8537
rect 3606 8463 3608 8472
rect 3660 8463 3662 8472
rect 3608 8434 3660 8440
rect 3606 7304 3662 7313
rect 3606 7239 3662 7248
rect 3514 6896 3570 6905
rect 3514 6831 3570 6840
rect 3528 5778 3556 6831
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3528 3738 3556 5510
rect 3620 4321 3648 7239
rect 3712 7206 3740 9998
rect 3804 9602 3832 12794
rect 3896 12306 3924 13087
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3882 12200 3938 12209
rect 3882 12135 3884 12144
rect 3936 12135 3938 12144
rect 3884 12106 3936 12112
rect 3882 10976 3938 10985
rect 3882 10911 3938 10920
rect 3896 10266 3924 10911
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3988 10112 4016 13670
rect 4080 13161 4108 14028
rect 4066 13152 4122 13161
rect 4066 13087 4122 13096
rect 4172 12986 4200 14758
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4068 12776 4120 12782
rect 4060 12724 4068 12764
rect 4060 12718 4120 12724
rect 4060 12702 4108 12718
rect 4080 12073 4108 12702
rect 4160 12436 4212 12442
rect 4264 12424 4292 20402
rect 4342 20360 4398 20369
rect 4342 20295 4398 20304
rect 4356 19854 4384 20295
rect 4344 19848 4396 19854
rect 4528 19848 4580 19854
rect 4344 19790 4396 19796
rect 4448 19808 4528 19836
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4356 17241 4384 19654
rect 4342 17232 4398 17241
rect 4342 17167 4398 17176
rect 4448 17082 4476 19808
rect 4528 19790 4580 19796
rect 4632 19666 4660 20538
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 5724 20256 5776 20262
rect 5816 20256 5868 20262
rect 5724 20198 5776 20204
rect 5814 20224 5816 20233
rect 5868 20224 5870 20233
rect 4710 20088 4766 20097
rect 4816 20058 4844 20198
rect 5538 20088 5594 20097
rect 4710 20023 4766 20032
rect 4804 20052 4856 20058
rect 4724 19689 4752 20023
rect 5538 20023 5594 20032
rect 4804 19994 4856 20000
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 4540 19638 4660 19666
rect 4710 19680 4766 19689
rect 4540 19514 4568 19638
rect 4710 19615 4766 19624
rect 4898 19612 5206 19621
rect 4898 19610 4904 19612
rect 4960 19610 4984 19612
rect 5040 19610 5064 19612
rect 5120 19610 5144 19612
rect 5200 19610 5206 19612
rect 4960 19558 4962 19610
rect 5142 19558 5144 19610
rect 4898 19556 4904 19558
rect 4960 19556 4984 19558
rect 5040 19556 5064 19558
rect 5120 19556 5144 19558
rect 5200 19556 5206 19558
rect 4898 19547 5206 19556
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4632 19468 5028 19496
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 4356 17054 4476 17082
rect 4356 15434 4384 17054
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4344 15428 4396 15434
rect 4344 15370 4396 15376
rect 4448 14600 4476 16934
rect 4540 16590 4568 18566
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4540 16425 4568 16526
rect 4632 16454 4660 19468
rect 4710 19408 4766 19417
rect 4710 19343 4766 19352
rect 4724 19281 4752 19343
rect 4710 19272 4766 19281
rect 4710 19207 4766 19216
rect 4804 19168 4856 19174
rect 5000 19156 5028 19468
rect 5264 19440 5316 19446
rect 5262 19408 5264 19417
rect 5316 19408 5318 19417
rect 5262 19343 5318 19352
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5172 19168 5224 19174
rect 5000 19128 5172 19156
rect 4804 19110 4856 19116
rect 5172 19110 5224 19116
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4724 18465 4752 18906
rect 4710 18456 4766 18465
rect 4710 18391 4766 18400
rect 4712 17604 4764 17610
rect 4712 17546 4764 17552
rect 4620 16448 4672 16454
rect 4526 16416 4582 16425
rect 4620 16390 4672 16396
rect 4526 16351 4582 16360
rect 4528 16176 4580 16182
rect 4528 16118 4580 16124
rect 4540 15162 4568 16118
rect 4632 15337 4660 16390
rect 4618 15328 4674 15337
rect 4618 15263 4674 15272
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4540 14657 4568 15098
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4356 14572 4476 14600
rect 4526 14648 4582 14657
rect 4526 14583 4582 14592
rect 4356 12617 4384 14572
rect 4632 14532 4660 15030
rect 4540 14504 4660 14532
rect 4434 14376 4490 14385
rect 4434 14311 4490 14320
rect 4448 12628 4476 14311
rect 4540 13433 4568 14504
rect 4724 13818 4752 17546
rect 4816 16561 4844 19110
rect 4898 18524 5206 18533
rect 4898 18522 4904 18524
rect 4960 18522 4984 18524
rect 5040 18522 5064 18524
rect 5120 18522 5144 18524
rect 5200 18522 5206 18524
rect 4960 18470 4962 18522
rect 5142 18470 5144 18522
rect 4898 18468 4904 18470
rect 4960 18468 4984 18470
rect 5040 18468 5064 18470
rect 5120 18468 5144 18470
rect 5200 18468 5206 18470
rect 4898 18459 5206 18468
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17649 5212 18022
rect 5170 17640 5226 17649
rect 5170 17575 5226 17584
rect 4898 17436 5206 17445
rect 4898 17434 4904 17436
rect 4960 17434 4984 17436
rect 5040 17434 5064 17436
rect 5120 17434 5144 17436
rect 5200 17434 5206 17436
rect 4960 17382 4962 17434
rect 5142 17382 5144 17434
rect 4898 17380 4904 17382
rect 4960 17380 4984 17382
rect 5040 17380 5064 17382
rect 5120 17380 5144 17382
rect 5200 17380 5206 17382
rect 4898 17371 5206 17380
rect 4802 16552 4858 16561
rect 4802 16487 4858 16496
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4816 14521 4844 16390
rect 4898 16348 5206 16357
rect 4898 16346 4904 16348
rect 4960 16346 4984 16348
rect 5040 16346 5064 16348
rect 5120 16346 5144 16348
rect 5200 16346 5206 16348
rect 4960 16294 4962 16346
rect 5142 16294 5144 16346
rect 4898 16292 4904 16294
rect 4960 16292 4984 16294
rect 5040 16292 5064 16294
rect 5120 16292 5144 16294
rect 5200 16292 5206 16294
rect 4898 16283 5206 16292
rect 5078 15872 5134 15881
rect 5078 15807 5134 15816
rect 5092 15366 5120 15807
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 4898 15260 5206 15269
rect 4898 15258 4904 15260
rect 4960 15258 4984 15260
rect 5040 15258 5064 15260
rect 5120 15258 5144 15260
rect 5200 15258 5206 15260
rect 4960 15206 4962 15258
rect 5142 15206 5144 15258
rect 4898 15204 4904 15206
rect 4960 15204 4984 15206
rect 5040 15204 5064 15206
rect 5120 15204 5144 15206
rect 5200 15204 5206 15206
rect 4898 15195 5206 15204
rect 4894 14920 4950 14929
rect 4894 14855 4950 14864
rect 4802 14512 4858 14521
rect 4802 14447 4858 14456
rect 4908 14260 4936 14855
rect 4632 13790 4752 13818
rect 4816 14232 4936 14260
rect 4526 13424 4582 13433
rect 4526 13359 4528 13368
rect 4580 13359 4582 13368
rect 4528 13330 4580 13336
rect 4526 13288 4582 13297
rect 4526 13223 4582 13232
rect 4540 12782 4568 13223
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4528 12640 4580 12646
rect 4342 12608 4398 12617
rect 4342 12543 4398 12552
rect 4448 12600 4528 12628
rect 4264 12396 4384 12424
rect 4160 12378 4212 12384
rect 4066 12064 4122 12073
rect 4066 11999 4122 12008
rect 4066 11792 4122 11801
rect 4066 11727 4068 11736
rect 4120 11727 4122 11736
rect 4068 11698 4120 11704
rect 4172 11529 4200 12378
rect 4250 12200 4306 12209
rect 4356 12186 4384 12396
rect 4448 12306 4476 12600
rect 4528 12582 4580 12588
rect 4526 12472 4582 12481
rect 4526 12407 4582 12416
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4306 12158 4384 12186
rect 4434 12200 4490 12209
rect 4250 12135 4306 12144
rect 4434 12135 4490 12144
rect 4158 11520 4214 11529
rect 4158 11455 4214 11464
rect 4066 11384 4122 11393
rect 4066 11319 4122 11328
rect 4080 11286 4108 11319
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 4250 11248 4306 11257
rect 4250 11183 4252 11192
rect 4304 11183 4306 11192
rect 4252 11154 4304 11160
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4068 10124 4120 10130
rect 3988 10084 4068 10112
rect 4068 10066 4120 10072
rect 4172 9926 4200 11018
rect 4264 10062 4292 11154
rect 4448 10713 4476 12135
rect 4434 10704 4490 10713
rect 4434 10639 4490 10648
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4066 9752 4122 9761
rect 4066 9687 4068 9696
rect 4120 9687 4122 9696
rect 4068 9658 4120 9664
rect 3804 9574 4016 9602
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3896 9058 3924 9454
rect 3804 9030 3924 9058
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3712 6361 3740 7142
rect 3698 6352 3754 6361
rect 3698 6287 3754 6296
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3712 5574 3740 6190
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3606 4312 3662 4321
rect 3606 4247 3662 4256
rect 3712 3992 3740 5102
rect 3804 4826 3832 9030
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3792 4616 3844 4622
rect 3790 4584 3792 4593
rect 3844 4584 3846 4593
rect 3790 4519 3846 4528
rect 3792 4004 3844 4010
rect 3712 3964 3792 3992
rect 3792 3946 3844 3952
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3896 3641 3924 8842
rect 3698 3632 3754 3641
rect 3698 3567 3754 3576
rect 3882 3632 3938 3641
rect 3882 3567 3938 3576
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 2872 3334 2924 3340
rect 3344 3352 3464 3380
rect 2884 3058 2912 3334
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2924 2748 3232 2757
rect 2924 2746 2930 2748
rect 2986 2746 3010 2748
rect 3066 2746 3090 2748
rect 3146 2746 3170 2748
rect 3226 2746 3232 2748
rect 2986 2694 2988 2746
rect 3168 2694 3170 2746
rect 2924 2692 2930 2694
rect 2986 2692 3010 2694
rect 3066 2692 3090 2694
rect 3146 2692 3170 2694
rect 3226 2692 3232 2694
rect 2924 2683 3232 2692
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 2870 2544 2926 2553
rect 2688 2508 2740 2514
rect 2870 2479 2926 2488
rect 2688 2450 2740 2456
rect 2884 2446 2912 2479
rect 2872 2440 2924 2446
rect 2502 2408 2558 2417
rect 3160 2417 3188 2586
rect 2872 2382 2924 2388
rect 3146 2408 3202 2417
rect 2502 2343 2558 2352
rect 3146 2343 3202 2352
rect 2688 1896 2740 1902
rect 2686 1864 2688 1873
rect 2740 1864 2742 1873
rect 2686 1799 2742 1808
rect 3344 1766 3372 3352
rect 3528 2774 3556 3470
rect 3712 3466 3740 3567
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3436 2746 3556 2774
rect 3436 2038 3464 2746
rect 3424 2032 3476 2038
rect 3424 1974 3476 1980
rect 3804 1834 3832 3470
rect 3988 2394 4016 9574
rect 4264 9466 4292 9998
rect 4342 9616 4398 9625
rect 4342 9551 4398 9560
rect 4080 9438 4292 9466
rect 4080 8537 4108 9438
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4066 8528 4122 8537
rect 4172 8514 4200 9318
rect 4356 8838 4384 9551
rect 4448 9042 4476 10639
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4434 8664 4490 8673
rect 4434 8599 4490 8608
rect 4342 8528 4398 8537
rect 4172 8486 4292 8514
rect 4066 8463 4122 8472
rect 4068 8424 4120 8430
rect 4066 8392 4068 8401
rect 4120 8392 4122 8401
rect 4066 8327 4122 8336
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4080 7206 4108 8026
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6225 4108 6598
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4068 5704 4120 5710
rect 4066 5672 4068 5681
rect 4120 5672 4122 5681
rect 4066 5607 4122 5616
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 4758 4108 5510
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4080 2854 4108 4558
rect 4172 3670 4200 7686
rect 4264 4826 4292 8486
rect 4342 8463 4398 8472
rect 4356 6866 4384 8463
rect 4448 8430 4476 8599
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4158 3360 4214 3369
rect 4158 3295 4214 3304
rect 4172 2922 4200 3295
rect 4160 2916 4212 2922
rect 4160 2858 4212 2864
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 4080 2582 4108 2790
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 4158 2408 4214 2417
rect 3988 2366 4108 2394
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3792 1828 3844 1834
rect 3792 1770 3844 1776
rect 2780 1760 2832 1766
rect 2780 1702 2832 1708
rect 3332 1760 3384 1766
rect 3332 1702 3384 1708
rect 2320 1352 2372 1358
rect 2320 1294 2372 1300
rect 2332 746 2360 1294
rect 2792 814 2820 1702
rect 2924 1660 3232 1669
rect 2924 1658 2930 1660
rect 2986 1658 3010 1660
rect 3066 1658 3090 1660
rect 3146 1658 3170 1660
rect 3226 1658 3232 1660
rect 2986 1606 2988 1658
rect 3168 1606 3170 1658
rect 2924 1604 2930 1606
rect 2986 1604 3010 1606
rect 3066 1604 3090 1606
rect 3146 1604 3170 1606
rect 3226 1604 3232 1606
rect 2924 1595 3232 1604
rect 3240 1488 3292 1494
rect 3240 1430 3292 1436
rect 3252 1358 3280 1430
rect 2964 1352 3016 1358
rect 2962 1320 2964 1329
rect 3240 1352 3292 1358
rect 3016 1320 3018 1329
rect 3240 1294 3292 1300
rect 2962 1255 3018 1264
rect 3148 1216 3200 1222
rect 3148 1158 3200 1164
rect 2780 808 2832 814
rect 2780 750 2832 756
rect 2320 740 2372 746
rect 2320 682 2372 688
rect 2228 264 2280 270
rect 2228 206 2280 212
rect 3160 202 3188 1158
rect 3252 338 3280 1294
rect 3988 542 4016 2246
rect 4080 1902 4108 2366
rect 4158 2343 4214 2352
rect 4172 2038 4200 2343
rect 4160 2032 4212 2038
rect 4160 1974 4212 1980
rect 4264 1970 4292 3538
rect 4252 1964 4304 1970
rect 4252 1906 4304 1912
rect 4068 1896 4120 1902
rect 4068 1838 4120 1844
rect 4252 1828 4304 1834
rect 4252 1770 4304 1776
rect 4066 1592 4122 1601
rect 4066 1527 4122 1536
rect 4080 1358 4108 1527
rect 4264 1426 4292 1770
rect 4356 1426 4384 6326
rect 4448 4146 4476 7958
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4434 3904 4490 3913
rect 4434 3839 4490 3848
rect 4448 3058 4476 3839
rect 4540 3602 4568 12407
rect 4632 10810 4660 13790
rect 4712 13728 4764 13734
rect 4710 13696 4712 13705
rect 4764 13696 4766 13705
rect 4710 13631 4766 13640
rect 4710 13016 4766 13025
rect 4710 12951 4712 12960
rect 4764 12951 4766 12960
rect 4712 12922 4764 12928
rect 4816 12866 4844 14232
rect 4898 14172 5206 14181
rect 4898 14170 4904 14172
rect 4960 14170 4984 14172
rect 5040 14170 5064 14172
rect 5120 14170 5144 14172
rect 5200 14170 5206 14172
rect 4960 14118 4962 14170
rect 5142 14118 5144 14170
rect 4898 14116 4904 14118
rect 4960 14116 4984 14118
rect 5040 14116 5064 14118
rect 5120 14116 5144 14118
rect 5200 14116 5206 14118
rect 4898 14107 5206 14116
rect 4894 13832 4950 13841
rect 4894 13767 4950 13776
rect 4908 13297 4936 13767
rect 4894 13288 4950 13297
rect 4894 13223 4950 13232
rect 4898 13084 5206 13093
rect 4898 13082 4904 13084
rect 4960 13082 4984 13084
rect 5040 13082 5064 13084
rect 5120 13082 5144 13084
rect 5200 13082 5206 13084
rect 4960 13030 4962 13082
rect 5142 13030 5144 13082
rect 4898 13028 4904 13030
rect 4960 13028 4984 13030
rect 5040 13028 5064 13030
rect 5120 13028 5144 13030
rect 5200 13028 5206 13030
rect 4898 13019 5206 13028
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4724 12838 4844 12866
rect 4724 11898 4752 12838
rect 4908 12753 4936 12922
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 4894 12744 4950 12753
rect 4894 12679 4950 12688
rect 4802 12472 4858 12481
rect 4802 12407 4858 12416
rect 4816 12238 4844 12407
rect 4986 12336 5042 12345
rect 4986 12271 4988 12280
rect 5040 12271 5042 12280
rect 4988 12242 5040 12248
rect 4804 12232 4856 12238
rect 5092 12209 5120 12854
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5184 12617 5212 12786
rect 5170 12608 5226 12617
rect 5170 12543 5226 12552
rect 4804 12174 4856 12180
rect 5078 12200 5134 12209
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4816 11778 4844 12174
rect 5078 12135 5134 12144
rect 4898 11996 5206 12005
rect 4898 11994 4904 11996
rect 4960 11994 4984 11996
rect 5040 11994 5064 11996
rect 5120 11994 5144 11996
rect 5200 11994 5206 11996
rect 4960 11942 4962 11994
rect 5142 11942 5144 11994
rect 4898 11940 4904 11942
rect 4960 11940 4984 11942
rect 5040 11940 5064 11942
rect 5120 11940 5144 11942
rect 5200 11940 5206 11942
rect 4898 11931 5206 11940
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4724 11750 4844 11778
rect 4724 10985 4752 11750
rect 5092 11529 5120 11834
rect 5170 11792 5226 11801
rect 5170 11727 5172 11736
rect 5224 11727 5226 11736
rect 5172 11698 5224 11704
rect 5184 11558 5212 11698
rect 5172 11552 5224 11558
rect 5078 11520 5134 11529
rect 5172 11494 5224 11500
rect 5078 11455 5134 11464
rect 4802 11384 4858 11393
rect 4802 11319 4858 11328
rect 4710 10976 4766 10985
rect 4710 10911 4766 10920
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4710 10568 4766 10577
rect 4710 10503 4766 10512
rect 4618 10296 4674 10305
rect 4618 10231 4674 10240
rect 4632 7750 4660 10231
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4632 3482 4660 6598
rect 4724 3924 4752 10503
rect 4816 9382 4844 11319
rect 4898 10908 5206 10917
rect 4898 10906 4904 10908
rect 4960 10906 4984 10908
rect 5040 10906 5064 10908
rect 5120 10906 5144 10908
rect 5200 10906 5206 10908
rect 4960 10854 4962 10906
rect 5142 10854 5144 10906
rect 4898 10852 4904 10854
rect 4960 10852 4984 10854
rect 5040 10852 5064 10854
rect 5120 10852 5144 10854
rect 5200 10852 5206 10854
rect 4898 10843 5206 10852
rect 5172 10600 5224 10606
rect 4894 10568 4950 10577
rect 5172 10542 5224 10548
rect 4894 10503 4950 10512
rect 5080 10532 5132 10538
rect 4908 10470 4936 10503
rect 5080 10474 5132 10480
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 5092 10130 5120 10474
rect 5184 10266 5212 10542
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4898 9820 5206 9829
rect 4898 9818 4904 9820
rect 4960 9818 4984 9820
rect 5040 9818 5064 9820
rect 5120 9818 5144 9820
rect 5200 9818 5206 9820
rect 4960 9766 4962 9818
rect 5142 9766 5144 9818
rect 4898 9764 4904 9766
rect 4960 9764 4984 9766
rect 5040 9764 5064 9766
rect 5120 9764 5144 9766
rect 5200 9764 5206 9766
rect 4898 9755 5206 9764
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4898 8732 5206 8741
rect 4898 8730 4904 8732
rect 4960 8730 4984 8732
rect 5040 8730 5064 8732
rect 5120 8730 5144 8732
rect 5200 8730 5206 8732
rect 4960 8678 4962 8730
rect 5142 8678 5144 8730
rect 4898 8676 4904 8678
rect 4960 8676 4984 8678
rect 5040 8676 5064 8678
rect 5120 8676 5144 8678
rect 5200 8676 5206 8678
rect 4898 8667 5206 8676
rect 5276 8616 5304 19246
rect 5368 15162 5396 19926
rect 5446 19816 5502 19825
rect 5446 19751 5502 19760
rect 5460 16833 5488 19751
rect 5552 19514 5580 20023
rect 5632 19780 5684 19786
rect 5632 19722 5684 19728
rect 5644 19689 5672 19722
rect 5630 19680 5686 19689
rect 5630 19615 5686 19624
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5736 18873 5764 20198
rect 5814 20159 5870 20168
rect 6090 19952 6146 19961
rect 6090 19887 6146 19896
rect 6460 19916 6512 19922
rect 5816 19848 5868 19854
rect 5868 19808 5948 19836
rect 5816 19790 5868 19796
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5828 19174 5856 19654
rect 5920 19553 5948 19808
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 5906 19544 5962 19553
rect 5906 19479 5962 19488
rect 5908 19236 5960 19242
rect 5908 19178 5960 19184
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5722 18864 5778 18873
rect 5722 18799 5778 18808
rect 5736 18766 5764 18799
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5828 18630 5856 19110
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5630 18184 5686 18193
rect 5630 18119 5686 18128
rect 5446 16824 5502 16833
rect 5446 16759 5502 16768
rect 5448 16720 5500 16726
rect 5448 16662 5500 16668
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5354 14512 5410 14521
rect 5354 14447 5410 14456
rect 5368 12986 5396 14447
rect 5460 13326 5488 16662
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5552 15502 5580 16390
rect 5644 15706 5672 18119
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5736 17066 5764 17818
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 13394 5580 15438
rect 5632 14884 5684 14890
rect 5632 14826 5684 14832
rect 5644 14550 5672 14826
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5630 13696 5686 13705
rect 5630 13631 5686 13640
rect 5644 13530 5672 13631
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5460 12918 5488 13126
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5446 12744 5502 12753
rect 5356 12708 5408 12714
rect 5446 12679 5502 12688
rect 5540 12708 5592 12714
rect 5356 12650 5408 12656
rect 5368 10606 5396 12650
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5184 8588 5304 8616
rect 5184 8498 5212 8588
rect 5368 8548 5396 10542
rect 5460 9586 5488 12679
rect 5540 12650 5592 12656
rect 5552 11014 5580 12650
rect 5644 11642 5672 13262
rect 5736 11762 5764 15846
rect 5828 14056 5856 17478
rect 5920 16182 5948 19178
rect 6012 17202 6040 19654
rect 6104 19446 6132 19887
rect 6460 19858 6512 19864
rect 6092 19440 6144 19446
rect 6092 19382 6144 19388
rect 6090 19000 6146 19009
rect 6090 18935 6146 18944
rect 6104 18834 6132 18935
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5908 16176 5960 16182
rect 5908 16118 5960 16124
rect 5908 15972 5960 15978
rect 5908 15914 5960 15920
rect 5920 15094 5948 15914
rect 5908 15088 5960 15094
rect 5908 15030 5960 15036
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5920 14414 5948 14758
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5828 14028 5948 14056
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5828 13433 5856 13874
rect 5814 13424 5870 13433
rect 5814 13359 5870 13368
rect 5920 13190 5948 14028
rect 5908 13184 5960 13190
rect 5814 13152 5870 13161
rect 5908 13126 5960 13132
rect 5814 13087 5870 13096
rect 5828 12850 5856 13087
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5828 11694 5856 12786
rect 5920 12102 5948 12922
rect 6012 12714 6040 16934
rect 6104 15366 6132 17682
rect 6196 16794 6224 18702
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6288 18329 6316 18362
rect 6472 18358 6500 19858
rect 6642 19816 6698 19825
rect 6642 19751 6698 19760
rect 6550 19408 6606 19417
rect 6656 19378 6684 19751
rect 6550 19343 6606 19352
rect 6644 19372 6696 19378
rect 6564 18850 6592 19343
rect 6644 19314 6696 19320
rect 6564 18822 6684 18850
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6460 18352 6512 18358
rect 6274 18320 6330 18329
rect 6460 18294 6512 18300
rect 6274 18255 6330 18264
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6288 17882 6316 18022
rect 6366 17912 6422 17921
rect 6276 17876 6328 17882
rect 6366 17847 6422 17856
rect 6276 17818 6328 17824
rect 6380 17513 6408 17847
rect 6472 17592 6500 18294
rect 6564 18057 6592 18702
rect 6550 18048 6606 18057
rect 6550 17983 6606 17992
rect 6552 17604 6604 17610
rect 6472 17564 6552 17592
rect 6552 17546 6604 17552
rect 6366 17504 6422 17513
rect 6366 17439 6422 17448
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6472 17241 6500 17274
rect 6458 17232 6514 17241
rect 6276 17196 6328 17202
rect 6458 17167 6514 17176
rect 6276 17138 6328 17144
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 6092 15360 6144 15366
rect 6092 15302 6144 15308
rect 6090 15192 6146 15201
rect 6090 15127 6146 15136
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5816 11688 5868 11694
rect 5644 11614 5764 11642
rect 5816 11630 5868 11636
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 8673 5488 9318
rect 5446 8664 5502 8673
rect 5446 8599 5502 8608
rect 5276 8520 5396 8548
rect 5448 8560 5500 8566
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5078 8392 5134 8401
rect 5078 8327 5080 8336
rect 5132 8327 5134 8336
rect 5080 8298 5132 8304
rect 5092 7886 5120 8298
rect 5080 7880 5132 7886
rect 4802 7848 4858 7857
rect 5080 7822 5132 7828
rect 4802 7783 4804 7792
rect 4856 7783 4858 7792
rect 4804 7754 4856 7760
rect 4898 7644 5206 7653
rect 4898 7642 4904 7644
rect 4960 7642 4984 7644
rect 5040 7642 5064 7644
rect 5120 7642 5144 7644
rect 5200 7642 5206 7644
rect 4960 7590 4962 7642
rect 5142 7590 5144 7642
rect 4898 7588 4904 7590
rect 4960 7588 4984 7590
rect 5040 7588 5064 7590
rect 5120 7588 5144 7590
rect 5200 7588 5206 7590
rect 4898 7579 5206 7588
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 5184 6798 5212 6870
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4816 4049 4844 6666
rect 4898 6556 5206 6565
rect 4898 6554 4904 6556
rect 4960 6554 4984 6556
rect 5040 6554 5064 6556
rect 5120 6554 5144 6556
rect 5200 6554 5206 6556
rect 4960 6502 4962 6554
rect 5142 6502 5144 6554
rect 4898 6500 4904 6502
rect 4960 6500 4984 6502
rect 5040 6500 5064 6502
rect 5120 6500 5144 6502
rect 5200 6500 5206 6502
rect 4898 6491 5206 6500
rect 4898 5468 5206 5477
rect 4898 5466 4904 5468
rect 4960 5466 4984 5468
rect 5040 5466 5064 5468
rect 5120 5466 5144 5468
rect 5200 5466 5206 5468
rect 4960 5414 4962 5466
rect 5142 5414 5144 5466
rect 4898 5412 4904 5414
rect 4960 5412 4984 5414
rect 5040 5412 5064 5414
rect 5120 5412 5144 5414
rect 5200 5412 5206 5414
rect 4898 5403 5206 5412
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 5092 4826 5120 5170
rect 5170 5128 5226 5137
rect 5170 5063 5226 5072
rect 5184 5030 5212 5063
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4898 4380 5206 4389
rect 4898 4378 4904 4380
rect 4960 4378 4984 4380
rect 5040 4378 5064 4380
rect 5120 4378 5144 4380
rect 5200 4378 5206 4380
rect 4960 4326 4962 4378
rect 5142 4326 5144 4378
rect 4898 4324 4904 4326
rect 4960 4324 4984 4326
rect 5040 4324 5064 4326
rect 5120 4324 5144 4326
rect 5200 4324 5206 4326
rect 4898 4315 5206 4324
rect 4802 4040 4858 4049
rect 4802 3975 4858 3984
rect 4724 3896 4844 3924
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4540 3454 4660 3482
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4434 2816 4490 2825
rect 4434 2751 4490 2760
rect 4448 2310 4476 2751
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4252 1420 4304 1426
rect 4252 1362 4304 1368
rect 4344 1420 4396 1426
rect 4344 1362 4396 1368
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 3976 536 4028 542
rect 3976 478 4028 484
rect 4448 474 4476 2246
rect 4540 1494 4568 3454
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4632 2310 4660 3130
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 4724 1494 4752 3606
rect 4816 2038 4844 3896
rect 4898 3292 5206 3301
rect 4898 3290 4904 3292
rect 4960 3290 4984 3292
rect 5040 3290 5064 3292
rect 5120 3290 5144 3292
rect 5200 3290 5206 3292
rect 4960 3238 4962 3290
rect 5142 3238 5144 3290
rect 4898 3236 4904 3238
rect 4960 3236 4984 3238
rect 5040 3236 5064 3238
rect 5120 3236 5144 3238
rect 5200 3236 5206 3238
rect 4898 3227 5206 3236
rect 5172 2848 5224 2854
rect 5276 2836 5304 8520
rect 5448 8502 5500 8508
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 6254 5396 7686
rect 5460 6798 5488 8502
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5368 5030 5396 6054
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5224 2808 5304 2836
rect 5172 2790 5224 2796
rect 4898 2204 5206 2213
rect 4898 2202 4904 2204
rect 4960 2202 4984 2204
rect 5040 2202 5064 2204
rect 5120 2202 5144 2204
rect 5200 2202 5206 2204
rect 4960 2150 4962 2202
rect 5142 2150 5144 2202
rect 4898 2148 4904 2150
rect 4960 2148 4984 2150
rect 5040 2148 5064 2150
rect 5120 2148 5144 2150
rect 5200 2148 5206 2150
rect 4898 2139 5206 2148
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 5172 1964 5224 1970
rect 5172 1906 5224 1912
rect 5080 1896 5132 1902
rect 5184 1873 5212 1906
rect 5080 1838 5132 1844
rect 5170 1864 5226 1873
rect 5092 1562 5120 1838
rect 5170 1799 5226 1808
rect 5080 1556 5132 1562
rect 5080 1498 5132 1504
rect 4528 1488 4580 1494
rect 4528 1430 4580 1436
rect 4712 1488 4764 1494
rect 4712 1430 4764 1436
rect 5172 1352 5224 1358
rect 5224 1300 5304 1306
rect 5172 1294 5304 1300
rect 5184 1278 5304 1294
rect 4620 1216 4672 1222
rect 4620 1158 4672 1164
rect 4632 882 4660 1158
rect 4898 1116 5206 1125
rect 4898 1114 4904 1116
rect 4960 1114 4984 1116
rect 5040 1114 5064 1116
rect 5120 1114 5144 1116
rect 5200 1114 5206 1116
rect 4960 1062 4962 1114
rect 5142 1062 5144 1114
rect 4898 1060 4904 1062
rect 4960 1060 4984 1062
rect 5040 1060 5064 1062
rect 5120 1060 5144 1062
rect 5200 1060 5206 1062
rect 4898 1051 5206 1060
rect 4620 876 4672 882
rect 4620 818 4672 824
rect 5276 746 5304 1278
rect 5368 1170 5396 4966
rect 5460 3534 5488 6734
rect 5552 6254 5580 10474
rect 5644 7449 5672 11494
rect 5736 10198 5764 11614
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5722 10024 5778 10033
rect 5722 9959 5778 9968
rect 5630 7440 5686 7449
rect 5630 7375 5686 7384
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5538 6080 5594 6089
rect 5538 6015 5594 6024
rect 5552 5710 5580 6015
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5538 5536 5594 5545
rect 5538 5471 5594 5480
rect 5552 4593 5580 5471
rect 5538 4584 5594 4593
rect 5538 4519 5594 4528
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5446 3224 5502 3233
rect 5446 3159 5502 3168
rect 5460 3126 5488 3159
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5460 1494 5488 2926
rect 5552 2922 5580 3946
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5644 2446 5672 7278
rect 5736 4010 5764 9959
rect 5828 9042 5856 11630
rect 5920 11286 5948 12038
rect 5998 11928 6054 11937
rect 5998 11863 6054 11872
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 6012 10305 6040 11863
rect 5998 10296 6054 10305
rect 5998 10231 6054 10240
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 5998 10160 6054 10169
rect 5920 9654 5948 10134
rect 5998 10095 6054 10104
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5920 6440 5948 9590
rect 6012 7410 6040 10095
rect 6104 9994 6132 15127
rect 6196 14958 6224 16050
rect 6288 15609 6316 17138
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6380 16454 6408 16594
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6274 15600 6330 15609
rect 6274 15535 6330 15544
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 6182 14648 6238 14657
rect 6182 14583 6238 14592
rect 6196 13025 6224 14583
rect 6182 13016 6238 13025
rect 6182 12951 6238 12960
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6196 12345 6224 12854
rect 6182 12336 6238 12345
rect 6182 12271 6238 12280
rect 6288 12186 6316 15030
rect 6380 13297 6408 15846
rect 6472 14929 6500 17070
rect 6564 15706 6592 17546
rect 6656 16998 6684 18822
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6656 16289 6684 16934
rect 6748 16425 6776 21830
rect 6872 21244 7180 21253
rect 6872 21242 6878 21244
rect 6934 21242 6958 21244
rect 7014 21242 7038 21244
rect 7094 21242 7118 21244
rect 7174 21242 7180 21244
rect 6934 21190 6936 21242
rect 7116 21190 7118 21242
rect 6872 21188 6878 21190
rect 6934 21188 6958 21190
rect 7014 21188 7038 21190
rect 7094 21188 7118 21190
rect 7174 21188 7180 21190
rect 6872 21179 7180 21188
rect 6872 20156 7180 20165
rect 6872 20154 6878 20156
rect 6934 20154 6958 20156
rect 7014 20154 7038 20156
rect 7094 20154 7118 20156
rect 7174 20154 7180 20156
rect 6934 20102 6936 20154
rect 7116 20102 7118 20154
rect 6872 20100 6878 20102
rect 6934 20100 6958 20102
rect 7014 20100 7038 20102
rect 7094 20100 7118 20102
rect 7174 20100 7180 20102
rect 6872 20091 7180 20100
rect 7472 19236 7524 19242
rect 7472 19178 7524 19184
rect 6872 19068 7180 19077
rect 6872 19066 6878 19068
rect 6934 19066 6958 19068
rect 7014 19066 7038 19068
rect 7094 19066 7118 19068
rect 7174 19066 7180 19068
rect 6934 19014 6936 19066
rect 7116 19014 7118 19066
rect 6872 19012 6878 19014
rect 6934 19012 6958 19014
rect 7014 19012 7038 19014
rect 7094 19012 7118 19014
rect 7174 19012 7180 19014
rect 6872 19003 7180 19012
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7116 18329 7144 18702
rect 7484 18426 7512 19178
rect 7654 18592 7710 18601
rect 7654 18527 7710 18536
rect 7472 18420 7524 18426
rect 7300 18380 7472 18408
rect 7102 18320 7158 18329
rect 7102 18255 7158 18264
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 6872 17980 7180 17989
rect 6872 17978 6878 17980
rect 6934 17978 6958 17980
rect 7014 17978 7038 17980
rect 7094 17978 7118 17980
rect 7174 17978 7180 17980
rect 6934 17926 6936 17978
rect 7116 17926 7118 17978
rect 6872 17924 6878 17926
rect 6934 17924 6958 17926
rect 7014 17924 7038 17926
rect 7094 17924 7118 17926
rect 7174 17924 7180 17926
rect 6872 17915 7180 17924
rect 7102 17640 7158 17649
rect 7102 17575 7104 17584
rect 7156 17575 7158 17584
rect 7104 17546 7156 17552
rect 6872 16892 7180 16901
rect 6872 16890 6878 16892
rect 6934 16890 6958 16892
rect 7014 16890 7038 16892
rect 7094 16890 7118 16892
rect 7174 16890 7180 16892
rect 6934 16838 6936 16890
rect 7116 16838 7118 16890
rect 6872 16836 6878 16838
rect 6934 16836 6958 16838
rect 7014 16836 7038 16838
rect 7094 16836 7118 16838
rect 7174 16836 7180 16838
rect 6872 16827 7180 16836
rect 6918 16688 6974 16697
rect 6918 16623 6974 16632
rect 6828 16448 6880 16454
rect 6734 16416 6790 16425
rect 6828 16390 6880 16396
rect 6734 16351 6790 16360
rect 6642 16280 6698 16289
rect 6642 16215 6698 16224
rect 6656 16114 6684 16215
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6656 15337 6684 15846
rect 6642 15328 6698 15337
rect 6642 15263 6698 15272
rect 6656 15144 6684 15263
rect 6564 15116 6684 15144
rect 6564 15026 6592 15116
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6458 14920 6514 14929
rect 6458 14855 6514 14864
rect 6656 14532 6684 14962
rect 6748 14657 6776 16050
rect 6840 15910 6868 16390
rect 6932 15910 6960 16623
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 7116 15978 7144 16458
rect 7208 16114 7236 18226
rect 7300 16454 7328 18380
rect 7472 18362 7524 18368
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7484 17746 7512 18158
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7392 17377 7420 17614
rect 7668 17513 7696 18527
rect 7930 18320 7986 18329
rect 7852 18278 7930 18306
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7654 17504 7710 17513
rect 7654 17439 7710 17448
rect 7378 17368 7434 17377
rect 7378 17303 7434 17312
rect 7656 17264 7708 17270
rect 7656 17206 7708 17212
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7392 16561 7420 17070
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7470 16824 7526 16833
rect 7470 16759 7526 16768
rect 7378 16552 7434 16561
rect 7378 16487 7434 16496
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7286 16280 7342 16289
rect 7286 16215 7342 16224
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6872 15804 7180 15813
rect 6872 15802 6878 15804
rect 6934 15802 6958 15804
rect 7014 15802 7038 15804
rect 7094 15802 7118 15804
rect 7174 15802 7180 15804
rect 6934 15750 6936 15802
rect 7116 15750 7118 15802
rect 6872 15748 6878 15750
rect 6934 15748 6958 15750
rect 7014 15748 7038 15750
rect 7094 15748 7118 15750
rect 7174 15748 7180 15750
rect 6872 15739 7180 15748
rect 7194 15056 7250 15065
rect 7194 14991 7196 15000
rect 7248 14991 7250 15000
rect 7196 14962 7248 14968
rect 6872 14716 7180 14725
rect 6872 14714 6878 14716
rect 6934 14714 6958 14716
rect 7014 14714 7038 14716
rect 7094 14714 7118 14716
rect 7174 14714 7180 14716
rect 6934 14662 6936 14714
rect 7116 14662 7118 14714
rect 6872 14660 6878 14662
rect 6934 14660 6958 14662
rect 7014 14660 7038 14662
rect 7094 14660 7118 14662
rect 7174 14660 7180 14662
rect 6734 14648 6790 14657
rect 6872 14651 7180 14660
rect 7300 14618 7328 16215
rect 6734 14583 6790 14592
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 6458 14512 6514 14521
rect 6656 14504 6776 14532
rect 6458 14447 6514 14456
rect 6472 14346 6500 14447
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6366 13288 6422 13297
rect 6366 13223 6422 13232
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6380 12889 6408 13126
rect 6366 12880 6422 12889
rect 6366 12815 6422 12824
rect 6366 12744 6422 12753
rect 6366 12679 6368 12688
rect 6420 12679 6422 12688
rect 6368 12650 6420 12656
rect 6196 12158 6316 12186
rect 6196 10538 6224 12158
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6288 11626 6316 12038
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6182 10432 6238 10441
rect 6182 10367 6238 10376
rect 6196 10198 6224 10367
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6092 9988 6144 9994
rect 6092 9930 6144 9936
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6104 9353 6132 9454
rect 6090 9344 6146 9353
rect 6090 9279 6146 9288
rect 6288 9178 6316 11222
rect 6380 9926 6408 12650
rect 6472 12345 6500 13874
rect 6564 12646 6592 14282
rect 6748 14249 6776 14504
rect 6734 14240 6790 14249
rect 6734 14175 6790 14184
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6656 13161 6684 14010
rect 6748 13512 6776 14175
rect 7024 13802 7052 14554
rect 7116 13938 7144 14554
rect 7392 14498 7420 16390
rect 7484 15065 7512 16759
rect 7470 15056 7526 15065
rect 7470 14991 7526 15000
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7484 14521 7512 14894
rect 7300 14470 7420 14498
rect 7470 14512 7526 14521
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 13938 7236 14214
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 6872 13628 7180 13637
rect 6872 13626 6878 13628
rect 6934 13626 6958 13628
rect 7014 13626 7038 13628
rect 7094 13626 7118 13628
rect 7174 13626 7180 13628
rect 6934 13574 6936 13626
rect 7116 13574 7118 13626
rect 6872 13572 6878 13574
rect 6934 13572 6958 13574
rect 7014 13572 7038 13574
rect 7094 13572 7118 13574
rect 7174 13572 7180 13574
rect 6872 13563 7180 13572
rect 7012 13524 7064 13530
rect 6748 13484 6868 13512
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6642 13152 6698 13161
rect 6642 13087 6698 13096
rect 6748 13002 6776 13262
rect 6656 12974 6776 13002
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6458 12336 6514 12345
rect 6458 12271 6514 12280
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6472 11286 6500 11698
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6104 8838 6132 9114
rect 6182 9072 6238 9081
rect 6182 9007 6238 9016
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5920 6412 6040 6440
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5828 4554 5856 6190
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5814 4448 5870 4457
rect 5814 4383 5870 4392
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5828 3890 5856 4383
rect 5736 3862 5856 3890
rect 5736 2990 5764 3862
rect 5814 3768 5870 3777
rect 5814 3703 5870 3712
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5828 2774 5856 3703
rect 5736 2746 5856 2774
rect 5736 2446 5764 2746
rect 5920 2582 5948 6258
rect 6012 3505 6040 6412
rect 6104 3942 6132 8230
rect 6196 8090 6224 9007
rect 6274 8936 6330 8945
rect 6274 8871 6330 8880
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6196 7993 6224 8026
rect 6182 7984 6238 7993
rect 6182 7919 6238 7928
rect 6182 7576 6238 7585
rect 6182 7511 6238 7520
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6196 3738 6224 7511
rect 6288 7342 6316 8871
rect 6380 8566 6408 9454
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6274 6624 6330 6633
rect 6274 6559 6330 6568
rect 6288 5302 6316 6559
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 5998 3496 6054 3505
rect 5998 3431 6054 3440
rect 5998 3088 6054 3097
rect 5998 3023 6054 3032
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5736 2088 5764 2382
rect 6012 2281 6040 3023
rect 5998 2272 6054 2281
rect 5998 2207 6054 2216
rect 6012 2106 6040 2207
rect 6104 2145 6132 3674
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6196 3097 6224 3402
rect 6182 3088 6238 3097
rect 6182 3023 6238 3032
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6090 2136 6146 2145
rect 5552 2060 5764 2088
rect 6000 2100 6052 2106
rect 5552 1970 5580 2060
rect 6090 2071 6146 2080
rect 6000 2042 6052 2048
rect 5540 1964 5592 1970
rect 5540 1906 5592 1912
rect 5448 1488 5500 1494
rect 5448 1430 5500 1436
rect 6000 1284 6052 1290
rect 5644 1244 6000 1272
rect 5644 1170 5672 1244
rect 6000 1226 6052 1232
rect 5368 1142 5672 1170
rect 6196 921 6224 2450
rect 6288 2038 6316 5238
rect 6380 4010 6408 8366
rect 6472 6730 6500 11018
rect 6564 9042 6592 12582
rect 6656 11801 6684 12974
rect 6840 12900 6868 13484
rect 7012 13466 7064 13472
rect 7024 13172 7052 13466
rect 7104 13184 7156 13190
rect 7024 13144 7104 13172
rect 7104 13126 7156 13132
rect 7010 13016 7066 13025
rect 7010 12951 7066 12960
rect 6748 12872 6868 12900
rect 6748 12434 6776 12872
rect 7024 12753 7052 12951
rect 7104 12776 7156 12782
rect 7010 12744 7066 12753
rect 7104 12718 7156 12724
rect 7010 12679 7066 12688
rect 7116 12628 7144 12718
rect 7208 12696 7236 13670
rect 7300 13530 7328 14470
rect 7470 14447 7526 14456
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7300 12986 7328 13330
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7392 12889 7420 14350
rect 7576 14074 7604 17002
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7484 13326 7512 13942
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7576 13172 7604 13466
rect 7484 13144 7604 13172
rect 7378 12880 7434 12889
rect 7378 12815 7434 12824
rect 7484 12782 7512 13144
rect 7564 12912 7616 12918
rect 7562 12880 7564 12889
rect 7616 12880 7618 12889
rect 7562 12815 7618 12824
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7208 12668 7420 12696
rect 7116 12600 7328 12628
rect 6872 12540 7180 12549
rect 6872 12538 6878 12540
rect 6934 12538 6958 12540
rect 7014 12538 7038 12540
rect 7094 12538 7118 12540
rect 7174 12538 7180 12540
rect 6934 12486 6936 12538
rect 7116 12486 7118 12538
rect 6872 12484 6878 12486
rect 6934 12484 6958 12486
rect 7014 12484 7038 12486
rect 7094 12484 7118 12486
rect 7174 12484 7180 12486
rect 6872 12475 7180 12484
rect 6748 12406 6868 12434
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6748 12209 6776 12242
rect 6734 12200 6790 12209
rect 6734 12135 6790 12144
rect 6840 12102 6868 12406
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6920 12232 6972 12238
rect 6918 12200 6920 12209
rect 6972 12200 6974 12209
rect 7024 12170 7052 12310
rect 6918 12135 6974 12144
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 6642 11792 6698 11801
rect 6642 11727 6698 11736
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6656 8906 6684 11727
rect 6872 11452 7180 11461
rect 6872 11450 6878 11452
rect 6934 11450 6958 11452
rect 7014 11450 7038 11452
rect 7094 11450 7118 11452
rect 7174 11450 7180 11452
rect 6934 11398 6936 11450
rect 7116 11398 7118 11450
rect 6872 11396 6878 11398
rect 6934 11396 6958 11398
rect 7014 11396 7038 11398
rect 7094 11396 7118 11398
rect 7174 11396 7180 11398
rect 6872 11387 7180 11396
rect 7102 11248 7158 11257
rect 7102 11183 7158 11192
rect 7116 11150 7144 11183
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6872 10364 7180 10373
rect 6872 10362 6878 10364
rect 6934 10362 6958 10364
rect 7014 10362 7038 10364
rect 7094 10362 7118 10364
rect 7174 10362 7180 10364
rect 6934 10310 6936 10362
rect 7116 10310 7118 10362
rect 6872 10308 6878 10310
rect 6934 10308 6958 10310
rect 7014 10308 7038 10310
rect 7094 10308 7118 10310
rect 7174 10308 7180 10310
rect 6872 10299 7180 10308
rect 7208 10062 7236 12038
rect 7300 11014 7328 12600
rect 7392 11393 7420 12668
rect 7470 12608 7526 12617
rect 7470 12543 7526 12552
rect 7484 11558 7512 12543
rect 7562 12336 7618 12345
rect 7562 12271 7618 12280
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7378 11384 7434 11393
rect 7378 11319 7434 11328
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 6748 8974 6776 9998
rect 6826 9752 6882 9761
rect 6826 9687 6882 9696
rect 6840 9382 6868 9687
rect 7300 9654 7328 10950
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6872 9276 7180 9285
rect 6872 9274 6878 9276
rect 6934 9274 6958 9276
rect 7014 9274 7038 9276
rect 7094 9274 7118 9276
rect 7174 9274 7180 9276
rect 6934 9222 6936 9274
rect 7116 9222 7118 9274
rect 6872 9220 6878 9222
rect 6934 9220 6958 9222
rect 7014 9220 7038 9222
rect 7094 9220 7118 9222
rect 7174 9220 7180 9222
rect 6872 9211 7180 9220
rect 7392 9092 7420 11154
rect 7300 9064 7420 9092
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 7104 8968 7156 8974
rect 7156 8928 7236 8956
rect 7104 8910 7156 8916
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 6734 8800 6790 8809
rect 6734 8735 6790 8744
rect 6550 7984 6606 7993
rect 6748 7970 6776 8735
rect 6872 8188 7180 8197
rect 6872 8186 6878 8188
rect 6934 8186 6958 8188
rect 7014 8186 7038 8188
rect 7094 8186 7118 8188
rect 7174 8186 7180 8188
rect 6934 8134 6936 8186
rect 7116 8134 7118 8186
rect 6872 8132 6878 8134
rect 6934 8132 6958 8134
rect 7014 8132 7038 8134
rect 7094 8132 7118 8134
rect 7174 8132 7180 8134
rect 6872 8123 7180 8132
rect 6550 7919 6606 7928
rect 6656 7942 6776 7970
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6460 6316 6512 6322
rect 6564 6304 6592 7919
rect 6512 6276 6592 6304
rect 6460 6258 6512 6264
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6564 5914 6592 6054
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6656 5778 6684 7942
rect 7010 7440 7066 7449
rect 7010 7375 7012 7384
rect 7064 7375 7066 7384
rect 7012 7346 7064 7352
rect 6872 7100 7180 7109
rect 6872 7098 6878 7100
rect 6934 7098 6958 7100
rect 7014 7098 7038 7100
rect 7094 7098 7118 7100
rect 7174 7098 7180 7100
rect 6934 7046 6936 7098
rect 7116 7046 7118 7098
rect 6872 7044 6878 7046
rect 6934 7044 6958 7046
rect 7014 7044 7038 7046
rect 7094 7044 7118 7046
rect 7174 7044 7180 7046
rect 6872 7035 7180 7044
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 5914 6776 6598
rect 7208 6497 7236 8928
rect 7300 7750 7328 9064
rect 7484 9024 7512 11222
rect 7392 8996 7512 9024
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7392 7562 7420 8996
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7484 7886 7512 8842
rect 7576 7886 7604 12271
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7392 7534 7512 7562
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7194 6488 7250 6497
rect 7194 6423 7250 6432
rect 7102 6352 7158 6361
rect 7102 6287 7104 6296
rect 7156 6287 7158 6296
rect 7196 6316 7248 6322
rect 7104 6258 7156 6264
rect 7196 6258 7248 6264
rect 6872 6012 7180 6021
rect 6872 6010 6878 6012
rect 6934 6010 6958 6012
rect 7014 6010 7038 6012
rect 7094 6010 7118 6012
rect 7174 6010 7180 6012
rect 6934 5958 6936 6010
rect 7116 5958 7118 6010
rect 6872 5956 6878 5958
rect 6934 5956 6958 5958
rect 7014 5956 7038 5958
rect 7094 5956 7118 5958
rect 7174 5956 7180 5958
rect 6872 5947 7180 5956
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6748 5409 6776 5850
rect 6458 5400 6514 5409
rect 6734 5400 6790 5409
rect 6458 5335 6460 5344
rect 6512 5335 6514 5344
rect 6552 5364 6604 5370
rect 6460 5306 6512 5312
rect 6734 5335 6790 5344
rect 7010 5400 7066 5409
rect 7010 5335 7066 5344
rect 6552 5306 6604 5312
rect 6564 5250 6592 5306
rect 7024 5302 7052 5335
rect 6472 5222 6592 5250
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 6472 4282 6500 5222
rect 6644 5160 6696 5166
rect 6642 5128 6644 5137
rect 6696 5128 6698 5137
rect 6828 5092 6880 5098
rect 6642 5063 6698 5072
rect 6748 5052 6828 5080
rect 6642 4720 6698 4729
rect 6642 4655 6698 4664
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 6458 3904 6514 3913
rect 6458 3839 6514 3848
rect 6472 3534 6500 3839
rect 6564 3602 6592 4490
rect 6656 3942 6684 4655
rect 6748 4486 6776 5052
rect 6828 5034 6880 5040
rect 6872 4924 7180 4933
rect 6872 4922 6878 4924
rect 6934 4922 6958 4924
rect 7014 4922 7038 4924
rect 7094 4922 7118 4924
rect 7174 4922 7180 4924
rect 6934 4870 6936 4922
rect 7116 4870 7118 4922
rect 6872 4868 6878 4870
rect 6934 4868 6958 4870
rect 7014 4868 7038 4870
rect 7094 4868 7118 4870
rect 7174 4868 7180 4870
rect 6872 4859 7180 4868
rect 6918 4720 6974 4729
rect 6918 4655 6974 4664
rect 6826 4584 6882 4593
rect 6826 4519 6882 4528
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6840 4078 6868 4519
rect 6932 4146 6960 4655
rect 7208 4146 7236 6258
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6644 3936 6696 3942
rect 6642 3904 6644 3913
rect 6696 3904 6698 3913
rect 6642 3839 6698 3848
rect 6872 3836 7180 3845
rect 6872 3834 6878 3836
rect 6934 3834 6958 3836
rect 7014 3834 7038 3836
rect 7094 3834 7118 3836
rect 7174 3834 7180 3836
rect 6934 3782 6936 3834
rect 7116 3782 7118 3834
rect 6872 3780 6878 3782
rect 6934 3780 6958 3782
rect 7014 3780 7038 3782
rect 7094 3780 7118 3782
rect 7174 3780 7180 3782
rect 6872 3771 7180 3780
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6550 3224 6606 3233
rect 6550 3159 6606 3168
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 6288 1601 6316 1974
rect 6274 1592 6330 1601
rect 6274 1527 6330 1536
rect 6460 1556 6512 1562
rect 6460 1498 6512 1504
rect 6368 1488 6420 1494
rect 6368 1430 6420 1436
rect 6182 912 6238 921
rect 6182 847 6238 856
rect 5264 740 5316 746
rect 5264 682 5316 688
rect 4436 468 4488 474
rect 4436 410 4488 416
rect 6380 406 6408 1430
rect 6472 1193 6500 1498
rect 6564 1290 6592 3159
rect 6656 3108 6684 3674
rect 7010 3360 7066 3369
rect 7010 3295 7066 3304
rect 7024 3194 7052 3295
rect 7116 3194 7144 3674
rect 7196 3664 7248 3670
rect 7300 3652 7328 7278
rect 7392 6322 7420 7414
rect 7484 7206 7512 7534
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7392 6089 7420 6122
rect 7378 6080 7434 6089
rect 7378 6015 7434 6024
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7392 4457 7420 5850
rect 7378 4448 7434 4457
rect 7378 4383 7434 4392
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7392 3913 7420 4082
rect 7378 3904 7434 3913
rect 7378 3839 7434 3848
rect 7248 3624 7328 3652
rect 7196 3606 7248 3612
rect 7288 3528 7340 3534
rect 7484 3482 7512 6938
rect 7576 6934 7604 7822
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7562 6488 7618 6497
rect 7668 6458 7696 17206
rect 7760 17134 7788 17614
rect 7852 17610 7880 18278
rect 8036 18290 8064 22034
rect 8576 21956 8628 21962
rect 8576 21898 8628 21904
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8312 18630 8340 18906
rect 8484 18896 8536 18902
rect 8482 18864 8484 18873
rect 8536 18864 8538 18873
rect 8482 18799 8538 18808
rect 8482 18728 8538 18737
rect 8482 18663 8538 18672
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18290 8340 18566
rect 8496 18306 8524 18663
rect 8588 18426 8616 21898
rect 8846 21788 9154 21797
rect 8846 21786 8852 21788
rect 8908 21786 8932 21788
rect 8988 21786 9012 21788
rect 9068 21786 9092 21788
rect 9148 21786 9154 21788
rect 8908 21734 8910 21786
rect 9090 21734 9092 21786
rect 8846 21732 8852 21734
rect 8908 21732 8932 21734
rect 8988 21732 9012 21734
rect 9068 21732 9092 21734
rect 9148 21732 9154 21734
rect 8846 21723 9154 21732
rect 12794 21788 13102 21797
rect 12794 21786 12800 21788
rect 12856 21786 12880 21788
rect 12936 21786 12960 21788
rect 13016 21786 13040 21788
rect 13096 21786 13102 21788
rect 12856 21734 12858 21786
rect 13038 21734 13040 21786
rect 12794 21732 12800 21734
rect 12856 21732 12880 21734
rect 12936 21732 12960 21734
rect 13016 21732 13040 21734
rect 13096 21732 13102 21734
rect 12794 21723 13102 21732
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 8846 20700 9154 20709
rect 8846 20698 8852 20700
rect 8908 20698 8932 20700
rect 8988 20698 9012 20700
rect 9068 20698 9092 20700
rect 9148 20698 9154 20700
rect 8908 20646 8910 20698
rect 9090 20646 9092 20698
rect 8846 20644 8852 20646
rect 8908 20644 8932 20646
rect 8988 20644 9012 20646
rect 9068 20644 9092 20646
rect 9148 20644 9154 20646
rect 8846 20635 9154 20644
rect 8666 19680 8722 19689
rect 8666 19615 8722 19624
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 7930 18255 7986 18264
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8300 18284 8352 18290
rect 8496 18278 8616 18306
rect 8300 18226 8352 18232
rect 7930 17912 7986 17921
rect 8036 17898 8064 18226
rect 8116 18080 8168 18086
rect 8114 18048 8116 18057
rect 8168 18048 8170 18057
rect 8114 17983 8170 17992
rect 7986 17870 8064 17898
rect 7930 17847 7986 17856
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 8392 17808 8444 17814
rect 8392 17750 8444 17756
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7932 17196 7984 17202
rect 8036 17184 8064 17750
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 8128 17490 8156 17614
rect 8206 17504 8262 17513
rect 8128 17462 8206 17490
rect 8206 17439 8262 17448
rect 8036 17156 8156 17184
rect 7932 17138 7984 17144
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7760 15881 7788 16730
rect 7852 16697 7880 17138
rect 7944 16833 7972 17138
rect 8024 17060 8076 17066
rect 8024 17002 8076 17008
rect 7930 16824 7986 16833
rect 8036 16794 8064 17002
rect 7930 16759 7986 16768
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 7838 16688 7894 16697
rect 7838 16623 7894 16632
rect 8022 16280 8078 16289
rect 8128 16266 8156 17156
rect 8220 16454 8248 17439
rect 8298 17368 8354 17377
rect 8298 17303 8354 17312
rect 8312 16794 8340 17303
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8300 16584 8352 16590
rect 8298 16552 8300 16561
rect 8352 16552 8354 16561
rect 8298 16487 8354 16496
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8128 16238 8248 16266
rect 8022 16215 8024 16224
rect 8076 16215 8078 16224
rect 8024 16186 8076 16192
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 7746 15872 7802 15881
rect 7746 15807 7802 15816
rect 7748 15632 7800 15638
rect 7748 15574 7800 15580
rect 7760 14618 7788 15574
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7760 13841 7788 13942
rect 7746 13832 7802 13841
rect 7746 13767 7802 13776
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7852 13394 7880 13466
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7746 13016 7802 13025
rect 7746 12951 7802 12960
rect 7840 12980 7892 12986
rect 7760 12850 7788 12951
rect 7840 12922 7892 12928
rect 7852 12850 7880 12922
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7944 12753 7972 16050
rect 8128 15194 8156 16050
rect 8036 15166 8156 15194
rect 7746 12744 7802 12753
rect 7930 12744 7986 12753
rect 7746 12679 7802 12688
rect 7840 12708 7892 12714
rect 7760 8974 7788 12679
rect 7930 12679 7986 12688
rect 7840 12650 7892 12656
rect 7852 11218 7880 12650
rect 8036 12617 8064 15166
rect 8128 15094 8156 15166
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 8220 14770 8248 16238
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8312 16114 8340 16186
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8312 15570 8340 15846
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 15162 8340 15506
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8128 14742 8248 14770
rect 8022 12608 8078 12617
rect 8022 12543 8078 12552
rect 8128 12458 8156 14742
rect 8312 14600 8340 14962
rect 8220 14572 8340 14600
rect 8220 13569 8248 14572
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8206 13560 8262 13569
rect 8206 13495 8262 13504
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 7944 12430 8156 12458
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7852 8090 7880 11018
rect 7944 10538 7972 12430
rect 8024 12232 8076 12238
rect 8220 12209 8248 13194
rect 8024 12174 8076 12180
rect 8206 12200 8262 12209
rect 7932 10532 7984 10538
rect 7932 10474 7984 10480
rect 7944 10062 7972 10474
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7930 9752 7986 9761
rect 7930 9687 7986 9696
rect 7944 9364 7972 9687
rect 8036 9466 8064 12174
rect 8116 12164 8168 12170
rect 8206 12135 8262 12144
rect 8116 12106 8168 12112
rect 8128 11830 8156 12106
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 8128 10266 8156 11766
rect 8220 11762 8248 12038
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8206 11384 8262 11393
rect 8206 11319 8262 11328
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8114 10024 8170 10033
rect 8114 9959 8170 9968
rect 8128 9654 8156 9959
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8036 9438 8156 9466
rect 7944 9336 8064 9364
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7852 7478 7880 8026
rect 7944 7750 7972 9114
rect 8036 7886 8064 9336
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7840 7472 7892 7478
rect 7932 7472 7984 7478
rect 7840 7414 7892 7420
rect 7930 7440 7932 7449
rect 7984 7440 7986 7449
rect 7748 7404 7800 7410
rect 7930 7375 7986 7384
rect 7748 7346 7800 7352
rect 7562 6423 7618 6432
rect 7656 6452 7708 6458
rect 7288 3470 7340 3476
rect 7300 3346 7328 3470
rect 7392 3466 7512 3482
rect 7380 3460 7512 3466
rect 7432 3454 7512 3460
rect 7380 3402 7432 3408
rect 7576 3398 7604 6423
rect 7656 6394 7708 6400
rect 7760 6338 7788 7346
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7668 6310 7788 6338
rect 7668 5574 7696 6310
rect 7852 5914 7880 6802
rect 7944 5914 7972 7210
rect 8022 7168 8078 7177
rect 8022 7103 8078 7112
rect 8036 6798 8064 7103
rect 8024 6792 8076 6798
rect 8128 6769 8156 9438
rect 8024 6734 8076 6740
rect 8114 6760 8170 6769
rect 8114 6695 8170 6704
rect 8220 6497 8248 11319
rect 8312 10305 8340 14418
rect 8404 11744 8432 17750
rect 8588 17746 8616 18278
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8576 17604 8628 17610
rect 8576 17546 8628 17552
rect 8496 16969 8524 17546
rect 8588 17513 8616 17546
rect 8574 17504 8630 17513
rect 8574 17439 8630 17448
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8482 16960 8538 16969
rect 8482 16895 8538 16904
rect 8588 16590 8616 17070
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8680 16522 8708 19615
rect 8846 19612 9154 19621
rect 8846 19610 8852 19612
rect 8908 19610 8932 19612
rect 8988 19610 9012 19612
rect 9068 19610 9092 19612
rect 9148 19610 9154 19612
rect 8908 19558 8910 19610
rect 9090 19558 9092 19610
rect 8846 19556 8852 19558
rect 8908 19556 8932 19558
rect 8988 19556 9012 19558
rect 9068 19556 9092 19558
rect 9148 19556 9154 19558
rect 8846 19547 9154 19556
rect 9218 19408 9274 19417
rect 9218 19343 9274 19352
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8772 18170 8800 18770
rect 8846 18524 9154 18533
rect 8846 18522 8852 18524
rect 8908 18522 8932 18524
rect 8988 18522 9012 18524
rect 9068 18522 9092 18524
rect 9148 18522 9154 18524
rect 8908 18470 8910 18522
rect 9090 18470 9092 18522
rect 8846 18468 8852 18470
rect 8908 18468 8932 18470
rect 8988 18468 9012 18470
rect 9068 18468 9092 18470
rect 9148 18468 9154 18470
rect 8846 18459 9154 18468
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 8772 18142 8892 18170
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8668 16516 8720 16522
rect 8668 16458 8720 16464
rect 8484 16448 8536 16454
rect 8536 16408 8616 16436
rect 8484 16390 8536 16396
rect 8482 16280 8538 16289
rect 8482 16215 8538 16224
rect 8496 16182 8524 16215
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8496 14929 8524 15438
rect 8482 14920 8538 14929
rect 8482 14855 8538 14864
rect 8588 14482 8616 16408
rect 8772 16402 8800 18022
rect 8864 17542 8892 18142
rect 9048 17610 9076 18362
rect 9232 17954 9260 19343
rect 9324 18426 9352 21354
rect 10820 21244 11128 21253
rect 10820 21242 10826 21244
rect 10882 21242 10906 21244
rect 10962 21242 10986 21244
rect 11042 21242 11066 21244
rect 11122 21242 11128 21244
rect 10882 21190 10884 21242
rect 11064 21190 11066 21242
rect 10820 21188 10826 21190
rect 10882 21188 10906 21190
rect 10962 21188 10986 21190
rect 11042 21188 11066 21190
rect 11122 21188 11128 21190
rect 10820 21179 11128 21188
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9508 18329 9536 18362
rect 9494 18320 9550 18329
rect 9494 18255 9550 18264
rect 9692 18057 9720 20402
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 9678 18048 9734 18057
rect 9678 17983 9734 17992
rect 9140 17926 9260 17954
rect 9140 17678 9168 17926
rect 9312 17876 9364 17882
rect 9508 17870 9812 17898
rect 9508 17864 9536 17870
rect 9364 17836 9536 17864
rect 9312 17818 9364 17824
rect 9588 17808 9640 17814
rect 9402 17776 9458 17785
rect 9220 17740 9272 17746
rect 9588 17750 9640 17756
rect 9402 17711 9458 17720
rect 9220 17682 9272 17688
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8846 17436 9154 17445
rect 8846 17434 8852 17436
rect 8908 17434 8932 17436
rect 8988 17434 9012 17436
rect 9068 17434 9092 17436
rect 9148 17434 9154 17436
rect 8908 17382 8910 17434
rect 9090 17382 9092 17434
rect 8846 17380 8852 17382
rect 8908 17380 8932 17382
rect 8988 17380 9012 17382
rect 9068 17380 9092 17382
rect 9148 17380 9154 17382
rect 8846 17371 9154 17380
rect 9232 17320 9260 17682
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9140 17292 9260 17320
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9048 17105 9076 17138
rect 9034 17096 9090 17105
rect 9034 17031 9090 17040
rect 8944 16720 8996 16726
rect 8944 16662 8996 16668
rect 8956 16590 8984 16662
rect 9140 16590 9168 17292
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 8680 16374 8800 16402
rect 8680 16096 8708 16374
rect 8846 16348 9154 16357
rect 8846 16346 8852 16348
rect 8908 16346 8932 16348
rect 8988 16346 9012 16348
rect 9068 16346 9092 16348
rect 9148 16346 9154 16348
rect 8908 16294 8910 16346
rect 9090 16294 9092 16346
rect 8846 16292 8852 16294
rect 8908 16292 8932 16294
rect 8988 16292 9012 16294
rect 9068 16292 9092 16294
rect 9148 16292 9154 16294
rect 8846 16283 9154 16292
rect 8760 16244 8812 16250
rect 8812 16204 8892 16232
rect 8760 16186 8812 16192
rect 8680 16068 8800 16096
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8680 15450 8708 15914
rect 8772 15910 8800 16068
rect 8864 15978 8892 16204
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 9034 15872 9090 15881
rect 9034 15807 9090 15816
rect 9048 15502 9076 15807
rect 9036 15496 9088 15502
rect 8942 15464 8998 15473
rect 8680 15422 8800 15450
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8496 13530 8524 14350
rect 8680 14346 8708 15302
rect 8772 14906 8800 15422
rect 9232 15473 9260 16458
rect 9324 16289 9352 17546
rect 9416 17066 9444 17711
rect 9600 17678 9628 17750
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9508 16969 9536 17546
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9692 17105 9720 17138
rect 9678 17096 9734 17105
rect 9678 17031 9734 17040
rect 9784 17048 9812 17870
rect 9862 17504 9918 17513
rect 9862 17439 9918 17448
rect 9876 17202 9904 17439
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9784 17020 9904 17048
rect 9680 16992 9732 16998
rect 9494 16960 9550 16969
rect 9494 16895 9550 16904
rect 9678 16960 9680 16969
rect 9732 16960 9734 16969
rect 9678 16895 9734 16904
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9310 16280 9366 16289
rect 9310 16215 9366 16224
rect 9404 16176 9456 16182
rect 9404 16118 9456 16124
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9324 15881 9352 15982
rect 9310 15872 9366 15881
rect 9310 15807 9366 15816
rect 9416 15502 9444 16118
rect 9508 15570 9536 16730
rect 9680 16448 9732 16454
rect 9678 16416 9680 16425
rect 9732 16416 9734 16425
rect 9678 16351 9734 16360
rect 9784 16250 9812 16730
rect 9876 16454 9904 17020
rect 9864 16448 9916 16454
rect 9968 16425 9996 18294
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10060 17377 10088 17478
rect 10046 17368 10102 17377
rect 10046 17303 10102 17312
rect 10046 17096 10102 17105
rect 10046 17031 10102 17040
rect 9864 16390 9916 16396
rect 9954 16416 10010 16425
rect 9954 16351 10010 16360
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9770 16144 9826 16153
rect 9588 16108 9640 16114
rect 9640 16068 9720 16096
rect 9770 16079 9826 16088
rect 9864 16108 9916 16114
rect 9588 16050 9640 16056
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9404 15496 9456 15502
rect 9036 15438 9088 15444
rect 9218 15464 9274 15473
rect 8942 15399 8998 15408
rect 9404 15438 9456 15444
rect 9494 15464 9550 15473
rect 9218 15399 9274 15408
rect 8956 15366 8984 15399
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 8846 15260 9154 15269
rect 8846 15258 8852 15260
rect 8908 15258 8932 15260
rect 8988 15258 9012 15260
rect 9068 15258 9092 15260
rect 9148 15258 9154 15260
rect 8908 15206 8910 15258
rect 9090 15206 9092 15258
rect 8846 15204 8852 15206
rect 8908 15204 8932 15206
rect 8988 15204 9012 15206
rect 9068 15204 9092 15206
rect 9148 15204 9154 15206
rect 8846 15195 9154 15204
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 8772 14878 8984 14906
rect 8956 14822 8984 14878
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8864 14618 8892 14758
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8760 14544 8812 14550
rect 8758 14512 8760 14521
rect 8812 14512 8814 14521
rect 8758 14447 8814 14456
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8668 14340 8720 14346
rect 8668 14282 8720 14288
rect 8588 14249 8616 14282
rect 8956 14260 8984 14758
rect 9048 14634 9076 15098
rect 9126 14784 9182 14793
rect 9232 14770 9260 15302
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9324 15026 9352 15098
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9310 14920 9366 14929
rect 9310 14855 9366 14864
rect 9182 14742 9260 14770
rect 9126 14719 9182 14728
rect 9048 14606 9168 14634
rect 9140 14550 9168 14606
rect 9036 14544 9088 14550
rect 9128 14544 9180 14550
rect 9036 14486 9088 14492
rect 9126 14512 9128 14521
rect 9180 14512 9182 14521
rect 9048 14414 9076 14486
rect 9126 14447 9182 14456
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 8574 14240 8630 14249
rect 8574 14175 8630 14184
rect 8772 14232 8984 14260
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8496 13025 8524 13194
rect 8482 13016 8538 13025
rect 8482 12951 8538 12960
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8496 12102 8524 12854
rect 8588 12288 8616 13670
rect 8680 13326 8708 13738
rect 8772 13326 8800 14232
rect 8846 14172 9154 14181
rect 8846 14170 8852 14172
rect 8908 14170 8932 14172
rect 8988 14170 9012 14172
rect 9068 14170 9092 14172
rect 9148 14170 9154 14172
rect 8908 14118 8910 14170
rect 9090 14118 9092 14170
rect 8846 14116 8852 14118
rect 8908 14116 8932 14118
rect 8988 14116 9012 14118
rect 9068 14116 9092 14118
rect 9148 14116 9154 14118
rect 8846 14107 9154 14116
rect 8944 14068 8996 14074
rect 8996 14028 9076 14056
rect 8944 14010 8996 14016
rect 8850 13832 8906 13841
rect 8850 13767 8906 13776
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8864 13172 8892 13767
rect 8942 13696 8998 13705
rect 8942 13631 8998 13640
rect 8956 13258 8984 13631
rect 9048 13258 9076 14028
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 9140 13569 9168 13942
rect 9126 13560 9182 13569
rect 9126 13495 9182 13504
rect 8944 13252 8996 13258
rect 8944 13194 8996 13200
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 8772 13144 8892 13172
rect 8666 13016 8722 13025
rect 8666 12951 8722 12960
rect 8680 12442 8708 12951
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8588 12260 8708 12288
rect 8574 12200 8630 12209
rect 8574 12135 8630 12144
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8404 11716 8524 11744
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8404 10713 8432 11562
rect 8496 10985 8524 11716
rect 8482 10976 8538 10985
rect 8482 10911 8538 10920
rect 8390 10704 8446 10713
rect 8390 10639 8446 10648
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8298 10296 8354 10305
rect 8298 10231 8354 10240
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8312 8498 8340 10134
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8298 8392 8354 8401
rect 8298 8327 8354 8336
rect 8312 8294 8340 8327
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8206 6488 8262 6497
rect 8206 6423 8262 6432
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7760 5766 8156 5794
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7564 3392 7616 3398
rect 7300 3318 7420 3346
rect 7564 3334 7616 3340
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 6736 3120 6788 3126
rect 6656 3080 6736 3108
rect 6736 3062 6788 3068
rect 6642 2544 6698 2553
rect 6748 2530 6776 3062
rect 7286 2816 7342 2825
rect 6872 2748 7180 2757
rect 7286 2751 7342 2760
rect 6872 2746 6878 2748
rect 6934 2746 6958 2748
rect 7014 2746 7038 2748
rect 7094 2746 7118 2748
rect 7174 2746 7180 2748
rect 6934 2694 6936 2746
rect 7116 2694 7118 2746
rect 6872 2692 6878 2694
rect 6934 2692 6958 2694
rect 7014 2692 7038 2694
rect 7094 2692 7118 2694
rect 7174 2692 7180 2694
rect 6872 2683 7180 2692
rect 7300 2530 7328 2751
rect 6698 2502 6776 2530
rect 6642 2479 6698 2488
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6656 1494 6684 2382
rect 6748 1970 6776 2502
rect 7024 2502 7328 2530
rect 7024 2038 7052 2502
rect 7392 2292 7420 3318
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7484 2446 7512 3062
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7576 2689 7604 2926
rect 7668 2774 7696 5510
rect 7760 3466 7788 5766
rect 8128 5710 8156 5766
rect 7932 5704 7984 5710
rect 8116 5704 8168 5710
rect 7984 5664 8064 5692
rect 7932 5646 7984 5652
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7852 4826 7880 5306
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7852 3058 7880 4762
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7668 2746 7788 2774
rect 7562 2680 7618 2689
rect 7562 2615 7618 2624
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7654 2408 7710 2417
rect 7576 2292 7604 2382
rect 7654 2343 7710 2352
rect 7392 2264 7604 2292
rect 7012 2032 7064 2038
rect 7012 1974 7064 1980
rect 6736 1964 6788 1970
rect 6736 1906 6788 1912
rect 7104 1828 7156 1834
rect 7156 1788 7328 1816
rect 7104 1770 7156 1776
rect 6872 1660 7180 1669
rect 6872 1658 6878 1660
rect 6934 1658 6958 1660
rect 7014 1658 7038 1660
rect 7094 1658 7118 1660
rect 7174 1658 7180 1660
rect 6934 1606 6936 1658
rect 7116 1606 7118 1658
rect 6872 1604 6878 1606
rect 6934 1604 6958 1606
rect 7014 1604 7038 1606
rect 7094 1604 7118 1606
rect 7174 1604 7180 1606
rect 6872 1595 7180 1604
rect 7300 1601 7328 1788
rect 7286 1592 7342 1601
rect 6736 1556 6788 1562
rect 6788 1516 7052 1544
rect 7286 1527 7342 1536
rect 6736 1498 6788 1504
rect 6644 1488 6696 1494
rect 7024 1465 7052 1516
rect 6644 1430 6696 1436
rect 6826 1456 6882 1465
rect 6826 1391 6882 1400
rect 7010 1456 7066 1465
rect 7010 1391 7066 1400
rect 6840 1358 6868 1391
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 6552 1284 6604 1290
rect 6552 1226 6604 1232
rect 6458 1184 6514 1193
rect 6458 1119 6514 1128
rect 6656 610 6684 1294
rect 7668 1222 7696 2343
rect 7656 1216 7708 1222
rect 7656 1158 7708 1164
rect 6644 604 6696 610
rect 6644 546 6696 552
rect 6368 400 6420 406
rect 6368 342 6420 348
rect 3240 332 3292 338
rect 3240 274 3292 280
rect 3148 196 3200 202
rect 3148 138 3200 144
rect 7760 66 7788 2746
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7852 1737 7880 2586
rect 7838 1728 7894 1737
rect 7838 1663 7894 1672
rect 7944 785 7972 5238
rect 8036 5137 8064 5664
rect 8116 5646 8168 5652
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8022 5128 8078 5137
rect 8022 5063 8078 5072
rect 8036 4690 8064 5063
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8036 4321 8064 4422
rect 8022 4312 8078 4321
rect 8022 4247 8078 4256
rect 8022 3768 8078 3777
rect 8022 3703 8078 3712
rect 8036 3670 8064 3703
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 8128 3534 8156 5510
rect 8220 4010 8248 6326
rect 8312 5545 8340 8230
rect 8404 7818 8432 10406
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8298 5536 8354 5545
rect 8298 5471 8354 5480
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8312 4593 8340 4694
rect 8298 4584 8354 4593
rect 8298 4519 8354 4528
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8312 3942 8340 4519
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8116 3528 8168 3534
rect 8022 3496 8078 3505
rect 8116 3470 8168 3476
rect 8022 3431 8078 3440
rect 8208 3460 8260 3466
rect 8036 3040 8064 3431
rect 8208 3402 8260 3408
rect 8220 3369 8248 3402
rect 8206 3360 8262 3369
rect 8206 3295 8262 3304
rect 8036 3012 8156 3040
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 8036 2650 8064 2858
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8128 1222 8156 3012
rect 8404 2938 8432 7142
rect 8496 5778 8524 10610
rect 8588 10470 8616 12135
rect 8680 11218 8708 12260
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8772 10674 8800 13144
rect 8846 13084 9154 13093
rect 8846 13082 8852 13084
rect 8908 13082 8932 13084
rect 8988 13082 9012 13084
rect 9068 13082 9092 13084
rect 9148 13082 9154 13084
rect 8908 13030 8910 13082
rect 9090 13030 9092 13082
rect 8846 13028 8852 13030
rect 8908 13028 8932 13030
rect 8988 13028 9012 13030
rect 9068 13028 9092 13030
rect 9148 13028 9154 13030
rect 8846 13019 9154 13028
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 9128 12980 9180 12986
rect 9232 12968 9260 14282
rect 9180 12940 9260 12968
rect 9128 12922 9180 12928
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8864 12646 8892 12786
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 9048 12209 9076 12922
rect 9220 12776 9272 12782
rect 9126 12744 9182 12753
rect 9220 12718 9272 12724
rect 9126 12679 9182 12688
rect 9034 12200 9090 12209
rect 9034 12135 9090 12144
rect 9140 12084 9168 12679
rect 9232 12481 9260 12718
rect 9324 12714 9352 14855
rect 9416 14278 9444 15438
rect 9494 15399 9550 15408
rect 9508 14278 9536 15399
rect 9404 14272 9456 14278
rect 9402 14240 9404 14249
rect 9496 14272 9548 14278
rect 9456 14240 9458 14249
rect 9496 14214 9548 14220
rect 9402 14175 9458 14184
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9218 12472 9274 12481
rect 9218 12407 9274 12416
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9140 12056 9260 12084
rect 8846 11996 9154 12005
rect 8846 11994 8852 11996
rect 8908 11994 8932 11996
rect 8988 11994 9012 11996
rect 9068 11994 9092 11996
rect 9148 11994 9154 11996
rect 8908 11942 8910 11994
rect 9090 11942 9092 11994
rect 8846 11940 8852 11942
rect 8908 11940 8932 11942
rect 8988 11940 9012 11942
rect 9068 11940 9092 11942
rect 9148 11940 9154 11942
rect 8846 11931 9154 11940
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9034 11112 9090 11121
rect 9034 11047 9036 11056
rect 9088 11047 9090 11056
rect 9036 11018 9088 11024
rect 9140 11014 9168 11698
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 8846 10908 9154 10917
rect 8846 10906 8852 10908
rect 8908 10906 8932 10908
rect 8988 10906 9012 10908
rect 9068 10906 9092 10908
rect 9148 10906 9154 10908
rect 8908 10854 8910 10906
rect 9090 10854 9092 10906
rect 8846 10852 8852 10854
rect 8908 10852 8932 10854
rect 8988 10852 9012 10854
rect 9068 10852 9092 10854
rect 9148 10852 9154 10854
rect 8846 10843 9154 10852
rect 9034 10704 9090 10713
rect 8760 10668 8812 10674
rect 9034 10639 9090 10648
rect 8760 10610 8812 10616
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 9048 10130 9076 10639
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8760 10056 8812 10062
rect 9232 10033 9260 12056
rect 9324 11257 9352 12378
rect 9416 12073 9444 13874
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9508 13161 9536 13806
rect 9494 13152 9550 13161
rect 9494 13087 9550 13096
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9508 12646 9536 12718
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9600 12345 9628 15846
rect 9692 15026 9720 16068
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 12374 9720 14758
rect 9784 14346 9812 16079
rect 9864 16050 9916 16056
rect 9876 15978 9904 16050
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9876 14940 9904 15302
rect 9968 15065 9996 15846
rect 10060 15502 10088 17031
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 9954 15056 10010 15065
rect 9954 14991 10010 15000
rect 9956 14952 10008 14958
rect 9876 14912 9956 14940
rect 9956 14894 10008 14900
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9876 13870 9904 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9968 13870 9996 14010
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9784 12918 9812 13738
rect 9864 13728 9916 13734
rect 9862 13696 9864 13705
rect 9916 13696 9918 13705
rect 9862 13631 9918 13640
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9876 13274 9904 13466
rect 9968 13394 9996 13466
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9876 13246 9996 13274
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9876 12918 9904 13126
rect 9968 13025 9996 13246
rect 9954 13016 10010 13025
rect 9954 12951 10010 12960
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9770 12744 9826 12753
rect 9770 12679 9826 12688
rect 9680 12368 9732 12374
rect 9586 12336 9642 12345
rect 9784 12345 9812 12679
rect 9680 12310 9732 12316
rect 9770 12336 9826 12345
rect 9586 12271 9642 12280
rect 9968 12288 9996 12786
rect 9770 12271 9826 12280
rect 9876 12260 9996 12288
rect 9680 12232 9732 12238
rect 9586 12200 9642 12209
rect 9508 12158 9586 12186
rect 9402 12064 9458 12073
rect 9402 11999 9458 12008
rect 9508 11880 9536 12158
rect 9680 12174 9732 12180
rect 9770 12200 9826 12209
rect 9586 12135 9642 12144
rect 9586 12064 9642 12073
rect 9586 11999 9642 12008
rect 9600 11898 9628 11999
rect 9499 11852 9536 11880
rect 9588 11892 9640 11898
rect 9499 11812 9527 11852
rect 9588 11834 9640 11840
rect 9416 11784 9527 11812
rect 9310 11248 9366 11257
rect 9310 11183 9366 11192
rect 9416 10962 9444 11784
rect 9600 11744 9628 11834
rect 9324 10934 9444 10962
rect 9508 11716 9628 11744
rect 9324 10266 9352 10934
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 8760 9998 8812 10004
rect 9218 10024 9274 10033
rect 8576 9920 8628 9926
rect 8574 9888 8576 9897
rect 8628 9888 8630 9897
rect 8574 9823 8630 9832
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8588 7721 8616 9114
rect 8680 8809 8708 9318
rect 8772 9081 8800 9998
rect 9218 9959 9274 9968
rect 8846 9820 9154 9829
rect 8846 9818 8852 9820
rect 8908 9818 8932 9820
rect 8988 9818 9012 9820
rect 9068 9818 9092 9820
rect 9148 9818 9154 9820
rect 8908 9766 8910 9818
rect 9090 9766 9092 9818
rect 8846 9764 8852 9766
rect 8908 9764 8932 9766
rect 8988 9764 9012 9766
rect 9068 9764 9092 9766
rect 9148 9764 9154 9766
rect 8846 9755 9154 9764
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8758 9072 8814 9081
rect 8864 9042 8892 9590
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 8758 9007 8814 9016
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 8666 8800 8722 8809
rect 8666 8735 8722 8744
rect 8846 8732 9154 8741
rect 8846 8730 8852 8732
rect 8908 8730 8932 8732
rect 8988 8730 9012 8732
rect 9068 8730 9092 8732
rect 9148 8730 9154 8732
rect 8908 8678 8910 8730
rect 9090 8678 9092 8730
rect 8846 8676 8852 8678
rect 8908 8676 8932 8678
rect 8988 8676 9012 8678
rect 9068 8676 9092 8678
rect 9148 8676 9154 8678
rect 8666 8664 8722 8673
rect 8846 8667 9154 8676
rect 8666 8599 8722 8608
rect 8680 7750 8708 8599
rect 8758 8256 8814 8265
rect 8758 8191 8814 8200
rect 9034 8256 9090 8265
rect 9034 8191 9090 8200
rect 8668 7744 8720 7750
rect 8574 7712 8630 7721
rect 8668 7686 8720 7692
rect 8574 7647 8630 7656
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8496 5409 8524 5578
rect 8482 5400 8538 5409
rect 8482 5335 8538 5344
rect 8496 4078 8524 5335
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8496 3505 8524 3878
rect 8482 3496 8538 3505
rect 8482 3431 8538 3440
rect 8404 2910 8524 2938
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8220 2553 8248 2586
rect 8300 2576 8352 2582
rect 8206 2544 8262 2553
rect 8300 2518 8352 2524
rect 8206 2479 8262 2488
rect 8206 2136 8262 2145
rect 8206 2071 8262 2080
rect 8116 1216 8168 1222
rect 8116 1158 8168 1164
rect 8220 785 8248 2071
rect 8312 1834 8340 2518
rect 8404 2281 8432 2790
rect 8390 2272 8446 2281
rect 8390 2207 8446 2216
rect 8300 1828 8352 1834
rect 8300 1770 8352 1776
rect 8496 1562 8524 2910
rect 8588 2038 8616 7142
rect 8680 7041 8708 7686
rect 8772 7460 8800 8191
rect 9048 7750 9076 8191
rect 9232 7993 9260 9046
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9324 8265 9352 8774
rect 9310 8256 9366 8265
rect 9310 8191 9366 8200
rect 9218 7984 9274 7993
rect 9416 7954 9444 9386
rect 9218 7919 9274 7928
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 8846 7644 9154 7653
rect 8846 7642 8852 7644
rect 8908 7642 8932 7644
rect 8988 7642 9012 7644
rect 9068 7642 9092 7644
rect 9148 7642 9154 7644
rect 8908 7590 8910 7642
rect 9090 7590 9092 7642
rect 8846 7588 8852 7590
rect 8908 7588 8932 7590
rect 8988 7588 9012 7590
rect 9068 7588 9092 7590
rect 9148 7588 9154 7590
rect 8846 7579 9154 7588
rect 8772 7432 8984 7460
rect 8956 7274 8984 7432
rect 8944 7268 8996 7274
rect 9232 7256 9260 7822
rect 9324 7426 9352 7822
rect 9508 7546 9536 11716
rect 9586 11248 9642 11257
rect 9586 11183 9642 11192
rect 9600 11082 9628 11183
rect 9692 11082 9720 12174
rect 9770 12135 9826 12144
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9784 11014 9812 12135
rect 9772 11008 9824 11014
rect 9678 10976 9734 10985
rect 9772 10950 9824 10956
rect 9678 10911 9734 10920
rect 9586 9752 9642 9761
rect 9586 9687 9588 9696
rect 9640 9687 9642 9696
rect 9588 9658 9640 9664
rect 9586 9208 9642 9217
rect 9586 9143 9642 9152
rect 9600 9042 9628 9143
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9586 8664 9642 8673
rect 9586 8599 9588 8608
rect 9640 8599 9642 8608
rect 9588 8570 9640 8576
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9324 7398 9536 7426
rect 8944 7210 8996 7216
rect 9048 7228 9260 7256
rect 8666 7032 8722 7041
rect 8666 6967 8722 6976
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8772 6458 8800 6938
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8864 6644 8892 6802
rect 8956 6798 8984 7210
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9048 6644 9076 7228
rect 9126 7168 9182 7177
rect 9126 7103 9182 7112
rect 9140 6730 9168 7103
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 8864 6616 9076 6644
rect 8846 6556 9154 6565
rect 8846 6554 8852 6556
rect 8908 6554 8932 6556
rect 8988 6554 9012 6556
rect 9068 6554 9092 6556
rect 9148 6554 9154 6556
rect 8908 6502 8910 6554
rect 9090 6502 9092 6554
rect 8846 6500 8852 6502
rect 8908 6500 8932 6502
rect 8988 6500 9012 6502
rect 9068 6500 9092 6502
rect 9148 6500 9154 6502
rect 8846 6491 9154 6500
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8666 6352 8722 6361
rect 9324 6322 9352 6734
rect 8666 6287 8722 6296
rect 9312 6316 9364 6322
rect 8680 5030 8708 6287
rect 9312 6258 9364 6264
rect 8944 6248 8996 6254
rect 9416 6225 9444 6802
rect 8944 6190 8996 6196
rect 9402 6216 9458 6225
rect 8850 5944 8906 5953
rect 8850 5879 8906 5888
rect 8864 5846 8892 5879
rect 8852 5840 8904 5846
rect 8956 5817 8984 6190
rect 9402 6151 9458 6160
rect 9508 6100 9536 7398
rect 9600 7206 9628 8366
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9588 6996 9640 7002
rect 9692 6984 9720 10911
rect 9770 10432 9826 10441
rect 9770 10367 9826 10376
rect 9784 7954 9812 10367
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9876 7857 9904 12260
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9968 11150 9996 12106
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9968 10198 9996 10610
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9862 7848 9918 7857
rect 9862 7783 9918 7792
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9876 7449 9904 7686
rect 9862 7440 9918 7449
rect 9862 7375 9918 7384
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9784 7177 9812 7210
rect 9770 7168 9826 7177
rect 9770 7103 9826 7112
rect 9640 6956 9720 6984
rect 9770 7032 9826 7041
rect 9770 6967 9826 6976
rect 9588 6938 9640 6944
rect 9588 6656 9640 6662
rect 9586 6624 9588 6633
rect 9640 6624 9642 6633
rect 9784 6610 9812 6967
rect 9968 6848 9996 9454
rect 10060 7041 10088 15302
rect 10152 12424 10180 17614
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10244 17338 10272 17478
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10336 16794 10364 17070
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10244 15008 10272 16118
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10336 15337 10364 15438
rect 10322 15328 10378 15337
rect 10322 15263 10378 15272
rect 10324 15020 10376 15026
rect 10244 14980 10324 15008
rect 10324 14962 10376 14968
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10244 12617 10272 13874
rect 10336 12850 10364 14962
rect 10428 14550 10456 20878
rect 12794 20700 13102 20709
rect 12794 20698 12800 20700
rect 12856 20698 12880 20700
rect 12936 20698 12960 20700
rect 13016 20698 13040 20700
rect 13096 20698 13102 20700
rect 12856 20646 12858 20698
rect 13038 20646 13040 20698
rect 12794 20644 12800 20646
rect 12856 20644 12880 20646
rect 12936 20644 12960 20646
rect 13016 20644 13040 20646
rect 13096 20644 13102 20646
rect 12794 20635 13102 20644
rect 10820 20156 11128 20165
rect 10820 20154 10826 20156
rect 10882 20154 10906 20156
rect 10962 20154 10986 20156
rect 11042 20154 11066 20156
rect 11122 20154 11128 20156
rect 10882 20102 10884 20154
rect 11064 20102 11066 20154
rect 10820 20100 10826 20102
rect 10882 20100 10906 20102
rect 10962 20100 10986 20102
rect 11042 20100 11066 20102
rect 11122 20100 11128 20102
rect 10820 20091 11128 20100
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10704 17882 10732 19314
rect 10820 19068 11128 19077
rect 10820 19066 10826 19068
rect 10882 19066 10906 19068
rect 10962 19066 10986 19068
rect 11042 19066 11066 19068
rect 11122 19066 11128 19068
rect 10882 19014 10884 19066
rect 11064 19014 11066 19066
rect 10820 19012 10826 19014
rect 10882 19012 10906 19014
rect 10962 19012 10986 19014
rect 11042 19012 11066 19014
rect 11122 19012 11128 19014
rect 10820 19003 11128 19012
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 12070 18592 12126 18601
rect 10796 18465 10824 18566
rect 12070 18527 12126 18536
rect 10782 18456 10838 18465
rect 10782 18391 10838 18400
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 10820 17980 11128 17989
rect 10820 17978 10826 17980
rect 10882 17978 10906 17980
rect 10962 17978 10986 17980
rect 11042 17978 11066 17980
rect 11122 17978 11128 17980
rect 10882 17926 10884 17978
rect 11064 17926 11066 17978
rect 10820 17924 10826 17926
rect 10882 17924 10906 17926
rect 10962 17924 10986 17926
rect 11042 17924 11066 17926
rect 11122 17924 11128 17926
rect 10820 17915 11128 17924
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 11518 17776 11574 17785
rect 11518 17711 11574 17720
rect 11150 17640 11206 17649
rect 11150 17575 11206 17584
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10600 16992 10652 16998
rect 10704 16969 10732 17274
rect 10600 16934 10652 16940
rect 10690 16960 10746 16969
rect 10520 16425 10548 16934
rect 10612 16833 10640 16934
rect 10690 16895 10746 16904
rect 10820 16892 11128 16901
rect 10820 16890 10826 16892
rect 10882 16890 10906 16892
rect 10962 16890 10986 16892
rect 11042 16890 11066 16892
rect 11122 16890 11128 16892
rect 10882 16838 10884 16890
rect 11064 16838 11066 16890
rect 10820 16836 10826 16838
rect 10882 16836 10906 16838
rect 10962 16836 10986 16838
rect 11042 16836 11066 16838
rect 11122 16836 11128 16838
rect 10598 16824 10654 16833
rect 10820 16827 11128 16836
rect 10598 16759 10654 16768
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10600 16652 10652 16658
rect 10796 16640 10824 16730
rect 10652 16612 10824 16640
rect 10600 16594 10652 16600
rect 10598 16552 10654 16561
rect 10598 16487 10654 16496
rect 10506 16416 10562 16425
rect 10506 16351 10562 16360
rect 10612 16250 10640 16487
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10612 16114 10640 16186
rect 10888 16114 10916 16390
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10612 15966 10824 15994
rect 10612 15881 10640 15966
rect 10796 15910 10824 15966
rect 10692 15904 10744 15910
rect 10598 15872 10654 15881
rect 10692 15846 10744 15852
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10598 15807 10654 15816
rect 10598 15736 10654 15745
rect 10598 15671 10654 15680
rect 10612 15434 10640 15671
rect 10600 15428 10652 15434
rect 10600 15370 10652 15376
rect 10506 15056 10562 15065
rect 10506 14991 10508 15000
rect 10560 14991 10562 15000
rect 10508 14962 10560 14968
rect 10600 14884 10652 14890
rect 10600 14826 10652 14832
rect 10506 14648 10562 14657
rect 10506 14583 10562 14592
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10520 14006 10548 14583
rect 10612 14550 10640 14826
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10704 14362 10732 15846
rect 10820 15804 11128 15813
rect 10820 15802 10826 15804
rect 10882 15802 10906 15804
rect 10962 15802 10986 15804
rect 11042 15802 11066 15804
rect 11122 15802 11128 15804
rect 10882 15750 10884 15802
rect 11064 15750 11066 15802
rect 10820 15748 10826 15750
rect 10882 15748 10906 15750
rect 10962 15748 10986 15750
rect 11042 15748 11066 15750
rect 11122 15748 11128 15750
rect 10820 15739 11128 15748
rect 10968 15632 11020 15638
rect 10782 15600 10838 15609
rect 10782 15535 10838 15544
rect 10966 15600 10968 15609
rect 11020 15600 11022 15609
rect 10966 15535 11022 15544
rect 11060 15564 11112 15570
rect 10796 15502 10824 15535
rect 11060 15506 11112 15512
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 11072 15201 11100 15506
rect 11058 15192 11114 15201
rect 11058 15127 11114 15136
rect 10820 14716 11128 14725
rect 10820 14714 10826 14716
rect 10882 14714 10906 14716
rect 10962 14714 10986 14716
rect 11042 14714 11066 14716
rect 11122 14714 11128 14716
rect 10882 14662 10884 14714
rect 11064 14662 11066 14714
rect 10820 14660 10826 14662
rect 10882 14660 10906 14662
rect 10962 14660 10986 14662
rect 11042 14660 11066 14662
rect 11122 14660 11128 14662
rect 10820 14651 11128 14660
rect 10782 14512 10838 14521
rect 10966 14512 11022 14521
rect 10876 14476 10928 14482
rect 10838 14456 10876 14464
rect 10782 14447 10876 14456
rect 10796 14436 10876 14447
rect 10966 14447 11022 14456
rect 10876 14418 10928 14424
rect 10612 14334 10732 14362
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10428 13394 10456 13806
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10324 12640 10376 12646
rect 10230 12608 10286 12617
rect 10324 12582 10376 12588
rect 10230 12543 10286 12552
rect 10152 12396 10272 12424
rect 10138 12336 10194 12345
rect 10138 12271 10194 12280
rect 10152 11286 10180 12271
rect 10244 12073 10272 12396
rect 10230 12064 10286 12073
rect 10230 11999 10286 12008
rect 10230 11928 10286 11937
rect 10336 11898 10364 12582
rect 10230 11863 10286 11872
rect 10324 11892 10376 11898
rect 10244 11558 10272 11863
rect 10324 11834 10376 11840
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10428 11370 10456 13126
rect 10612 12968 10640 14334
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10520 12940 10640 12968
rect 10520 12152 10548 12940
rect 10704 12850 10732 14214
rect 10980 13734 11008 14447
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10968 13728 11020 13734
rect 11072 13716 11100 14010
rect 11164 13818 11192 17575
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11256 14346 11284 15982
rect 11532 15910 11560 17711
rect 11702 16688 11758 16697
rect 11702 16623 11758 16632
rect 11716 16590 11744 16623
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11702 16280 11758 16289
rect 11702 16215 11758 16224
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11336 15904 11388 15910
rect 11520 15904 11572 15910
rect 11336 15846 11388 15852
rect 11518 15872 11520 15881
rect 11572 15872 11574 15881
rect 11348 15638 11376 15846
rect 11518 15807 11574 15816
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11440 15348 11468 15438
rect 11520 15360 11572 15366
rect 11440 15320 11520 15348
rect 11520 15302 11572 15308
rect 11348 15162 11560 15178
rect 11336 15156 11560 15162
rect 11388 15150 11560 15156
rect 11336 15098 11388 15104
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11440 14414 11468 15030
rect 11532 14618 11560 15150
rect 11624 15065 11652 16050
rect 11716 15910 11744 16215
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11702 15736 11758 15745
rect 11702 15671 11758 15680
rect 11716 15502 11744 15671
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11716 15162 11744 15302
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11610 15056 11666 15065
rect 11610 14991 11666 15000
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11348 13870 11376 14214
rect 11336 13864 11388 13870
rect 11164 13790 11284 13818
rect 11336 13806 11388 13812
rect 11072 13688 11192 13716
rect 10968 13670 11020 13676
rect 10820 13628 11128 13637
rect 10820 13626 10826 13628
rect 10882 13626 10906 13628
rect 10962 13626 10986 13628
rect 11042 13626 11066 13628
rect 11122 13626 11128 13628
rect 10882 13574 10884 13626
rect 11064 13574 11066 13626
rect 10820 13572 10826 13574
rect 10882 13572 10906 13574
rect 10962 13572 10986 13574
rect 11042 13572 11066 13574
rect 11122 13572 11128 13574
rect 10820 13563 11128 13572
rect 11164 13326 11192 13688
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10612 12356 10640 12786
rect 10796 12628 10824 13194
rect 10888 12782 10916 13262
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10980 12850 11008 13126
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10704 12600 10824 12628
rect 10704 12424 10732 12600
rect 10820 12540 11128 12549
rect 10820 12538 10826 12540
rect 10882 12538 10906 12540
rect 10962 12538 10986 12540
rect 11042 12538 11066 12540
rect 11122 12538 11128 12540
rect 10882 12486 10884 12538
rect 11064 12486 11066 12538
rect 10820 12484 10826 12486
rect 10882 12484 10906 12486
rect 10962 12484 10986 12486
rect 11042 12484 11066 12486
rect 11122 12484 11128 12486
rect 10820 12475 11128 12484
rect 10704 12396 11100 12424
rect 10612 12328 10824 12356
rect 11072 12345 11100 12396
rect 10520 12124 10732 12152
rect 10598 12064 10654 12073
rect 10598 11999 10654 12008
rect 10612 11898 10640 11999
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10244 11342 10456 11370
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10138 10704 10194 10713
rect 10138 10639 10140 10648
rect 10192 10639 10194 10648
rect 10140 10610 10192 10616
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10046 7032 10102 7041
rect 10046 6967 10102 6976
rect 9968 6820 10088 6848
rect 9954 6760 10010 6769
rect 9954 6695 10010 6704
rect 9784 6582 9904 6610
rect 9586 6559 9642 6568
rect 9876 6372 9904 6582
rect 9968 6497 9996 6695
rect 10060 6662 10088 6820
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9954 6488 10010 6497
rect 9954 6423 10010 6432
rect 9876 6344 9996 6372
rect 9416 6072 9536 6100
rect 9218 5944 9274 5953
rect 9218 5879 9274 5888
rect 8852 5782 8904 5788
rect 8942 5808 8998 5817
rect 8942 5743 8998 5752
rect 9232 5710 9260 5879
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9310 5672 9366 5681
rect 9310 5607 9312 5616
rect 9364 5607 9366 5616
rect 9312 5578 9364 5584
rect 9036 5568 9088 5574
rect 9088 5528 9260 5556
rect 9036 5510 9088 5516
rect 8846 5468 9154 5477
rect 8846 5466 8852 5468
rect 8908 5466 8932 5468
rect 8988 5466 9012 5468
rect 9068 5466 9092 5468
rect 9148 5466 9154 5468
rect 8908 5414 8910 5466
rect 9090 5414 9092 5466
rect 8846 5412 8852 5414
rect 8908 5412 8932 5414
rect 8988 5412 9012 5414
rect 9068 5412 9092 5414
rect 9148 5412 9154 5414
rect 8846 5403 9154 5412
rect 9128 5228 9180 5234
rect 9232 5216 9260 5528
rect 9232 5188 9352 5216
rect 9128 5170 9180 5176
rect 8758 5128 8814 5137
rect 8758 5063 8814 5072
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8680 4214 8708 4626
rect 8668 4208 8720 4214
rect 8668 4150 8720 4156
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8680 2990 8708 4014
rect 8772 3126 8800 5063
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8850 4856 8906 4865
rect 8850 4791 8906 4800
rect 8864 4486 8892 4791
rect 8956 4758 8984 4966
rect 9140 4758 9168 5170
rect 8944 4752 8996 4758
rect 8944 4694 8996 4700
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9140 4486 9168 4558
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 8846 4380 9154 4389
rect 8846 4378 8852 4380
rect 8908 4378 8932 4380
rect 8988 4378 9012 4380
rect 9068 4378 9092 4380
rect 9148 4378 9154 4380
rect 8908 4326 8910 4378
rect 9090 4326 9092 4378
rect 8846 4324 8852 4326
rect 8908 4324 8932 4326
rect 8988 4324 9012 4326
rect 9068 4324 9092 4326
rect 9148 4324 9154 4326
rect 8846 4315 9154 4324
rect 9324 4321 9352 5188
rect 9310 4312 9366 4321
rect 9310 4247 9366 4256
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8864 3942 8892 4082
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8956 3602 8984 4150
rect 9220 4140 9272 4146
rect 9416 4128 9444 6072
rect 9770 5944 9826 5953
rect 9600 5902 9770 5930
rect 9494 5264 9550 5273
rect 9494 5199 9550 5208
rect 9508 4690 9536 5199
rect 9600 5137 9628 5902
rect 9770 5879 9826 5888
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9586 5128 9642 5137
rect 9586 5063 9642 5072
rect 9692 4978 9720 5782
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9784 5273 9812 5646
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9968 5522 9996 6344
rect 10152 5522 10180 10406
rect 10244 5930 10272 11342
rect 10324 11280 10376 11286
rect 10324 11222 10376 11228
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10336 10044 10364 11222
rect 10428 10112 10456 11222
rect 10520 10470 10548 11834
rect 10704 11506 10732 12124
rect 10796 11898 10824 12328
rect 11058 12336 11114 12345
rect 10876 12300 10928 12306
rect 11058 12271 11114 12280
rect 10876 12242 10928 12248
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10888 11665 10916 12242
rect 11164 12220 11192 13262
rect 10980 12192 11192 12220
rect 10980 11937 11008 12192
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10966 11928 11022 11937
rect 10966 11863 11022 11872
rect 11072 11665 11100 12038
rect 10874 11656 10930 11665
rect 10874 11591 10930 11600
rect 11058 11656 11114 11665
rect 11058 11591 11114 11600
rect 10612 11478 10732 11506
rect 10612 11286 10640 11478
rect 10820 11452 11128 11461
rect 10820 11450 10826 11452
rect 10882 11450 10906 11452
rect 10962 11450 10986 11452
rect 11042 11450 11066 11452
rect 11122 11450 11128 11452
rect 10882 11398 10884 11450
rect 11064 11398 11066 11450
rect 10820 11396 10826 11398
rect 10882 11396 10906 11398
rect 10962 11396 10986 11398
rect 11042 11396 11066 11398
rect 11122 11396 11128 11398
rect 10820 11387 11128 11396
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10600 11280 10652 11286
rect 10600 11222 10652 11228
rect 10692 11144 10744 11150
rect 10598 11112 10654 11121
rect 10692 11086 10744 11092
rect 10598 11047 10654 11056
rect 10612 11014 10640 11047
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10598 10840 10654 10849
rect 10598 10775 10654 10784
rect 10612 10606 10640 10775
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10428 10084 10640 10112
rect 10336 10016 10456 10044
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10336 6780 10364 9658
rect 10428 9092 10456 10016
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 10520 9382 10548 9930
rect 10612 9722 10640 10084
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10704 9568 10732 11086
rect 10796 10470 10824 11290
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10888 10554 10916 11018
rect 10966 10976 11022 10985
rect 10966 10911 11022 10920
rect 10980 10810 11008 10911
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11164 10674 11192 12038
rect 11256 11082 11284 13790
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11334 13560 11390 13569
rect 11334 13495 11336 13504
rect 11388 13495 11390 13504
rect 11336 13466 11388 13472
rect 11440 13240 11468 13670
rect 11348 13212 11468 13240
rect 11348 13025 11376 13212
rect 11426 13152 11482 13161
rect 11426 13087 11482 13096
rect 11334 13016 11390 13025
rect 11334 12951 11390 12960
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11348 12442 11376 12786
rect 11440 12696 11468 13087
rect 11532 13025 11560 14282
rect 11624 14278 11652 14758
rect 11716 14278 11744 14894
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11808 14226 11836 18158
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11900 14521 11928 16050
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11886 14512 11942 14521
rect 11886 14447 11942 14456
rect 11808 14198 11928 14226
rect 11610 14104 11666 14113
rect 11794 14104 11850 14113
rect 11610 14039 11666 14048
rect 11716 14062 11794 14090
rect 11624 13326 11652 14039
rect 11716 13802 11744 14062
rect 11794 14039 11850 14048
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11612 13320 11664 13326
rect 11664 13280 11744 13308
rect 11612 13262 11664 13268
rect 11518 13016 11574 13025
rect 11518 12951 11574 12960
rect 11440 12668 11652 12696
rect 11518 12608 11574 12617
rect 11518 12543 11574 12552
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 10888 10526 11192 10554
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10820 10364 11128 10373
rect 10820 10362 10826 10364
rect 10882 10362 10906 10364
rect 10962 10362 10986 10364
rect 11042 10362 11066 10364
rect 11122 10362 11128 10364
rect 10882 10310 10884 10362
rect 11064 10310 11066 10362
rect 10820 10308 10826 10310
rect 10882 10308 10906 10310
rect 10962 10308 10986 10310
rect 11042 10308 11066 10310
rect 11122 10308 11128 10310
rect 10820 10299 11128 10308
rect 10704 9540 11008 9568
rect 10980 9518 11008 9540
rect 10980 9512 11036 9518
rect 10690 9480 10746 9489
rect 10980 9472 10984 9512
rect 10984 9454 11036 9460
rect 10690 9415 10746 9424
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 9110 10640 9318
rect 10600 9104 10652 9110
rect 10428 9064 10548 9092
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10428 7818 10456 8434
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10428 6882 10456 7754
rect 10520 7290 10548 9064
rect 10600 9046 10652 9052
rect 10704 8956 10732 9415
rect 10820 9276 11128 9285
rect 10820 9274 10826 9276
rect 10882 9274 10906 9276
rect 10962 9274 10986 9276
rect 11042 9274 11066 9276
rect 11122 9274 11128 9276
rect 10882 9222 10884 9274
rect 11064 9222 11066 9274
rect 10820 9220 10826 9222
rect 10882 9220 10906 9222
rect 10962 9220 10986 9222
rect 11042 9220 11066 9222
rect 11122 9220 11128 9222
rect 10820 9211 11128 9220
rect 11164 9042 11192 10526
rect 11244 10532 11296 10538
rect 11244 10474 11296 10480
rect 11256 10305 11284 10474
rect 11348 10441 11376 11834
rect 11440 11257 11468 11834
rect 11532 11642 11560 12543
rect 11624 11762 11652 12668
rect 11716 11937 11744 13280
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11808 12714 11836 13194
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 11794 12472 11850 12481
rect 11794 12407 11850 12416
rect 11702 11928 11758 11937
rect 11702 11863 11758 11872
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11532 11614 11652 11642
rect 11426 11248 11482 11257
rect 11426 11183 11482 11192
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11334 10432 11390 10441
rect 11334 10367 11390 10376
rect 11242 10296 11298 10305
rect 11242 10231 11298 10240
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11348 9722 11376 10202
rect 11440 10062 11468 11018
rect 11532 10606 11560 11086
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11532 10266 11560 10542
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 10612 8928 10732 8956
rect 10612 8004 10640 8928
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8276 10824 8774
rect 10874 8664 10930 8673
rect 10874 8599 10930 8608
rect 10888 8566 10916 8599
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10704 8248 10824 8276
rect 10704 8072 10732 8248
rect 10820 8188 11128 8197
rect 10820 8186 10826 8188
rect 10882 8186 10906 8188
rect 10962 8186 10986 8188
rect 11042 8186 11066 8188
rect 11122 8186 11128 8188
rect 10882 8134 10884 8186
rect 11064 8134 11066 8186
rect 10820 8132 10826 8134
rect 10882 8132 10906 8134
rect 10962 8132 10986 8134
rect 11042 8132 11066 8134
rect 11122 8132 11128 8134
rect 10820 8123 11128 8132
rect 10784 8084 10836 8090
rect 10704 8044 10784 8072
rect 10784 8026 10836 8032
rect 10612 7976 10732 8004
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10612 7410 10640 7754
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10520 7262 10640 7290
rect 10704 7274 10732 7976
rect 10782 7984 10838 7993
rect 10782 7919 10838 7928
rect 10796 7818 10824 7919
rect 10966 7848 11022 7857
rect 10784 7812 10836 7818
rect 10966 7783 11022 7792
rect 10784 7754 10836 7760
rect 10980 7449 11008 7783
rect 10966 7440 11022 7449
rect 10966 7375 11022 7384
rect 10428 6854 10548 6882
rect 10304 6752 10364 6780
rect 10304 6440 10332 6752
rect 10416 6452 10468 6458
rect 10304 6412 10364 6440
rect 10336 6254 10364 6412
rect 10416 6394 10468 6400
rect 10324 6248 10376 6254
rect 10428 6225 10456 6394
rect 10324 6190 10376 6196
rect 10414 6216 10470 6225
rect 10414 6151 10470 6160
rect 10324 6112 10376 6118
rect 10322 6080 10324 6089
rect 10520 6100 10548 6854
rect 10376 6080 10378 6089
rect 10322 6015 10378 6024
rect 10428 6072 10548 6100
rect 10244 5902 10364 5930
rect 10232 5840 10284 5846
rect 10230 5808 10232 5817
rect 10284 5808 10286 5817
rect 10230 5743 10286 5752
rect 9876 5302 9904 5510
rect 9968 5494 10088 5522
rect 10152 5494 10272 5522
rect 9864 5296 9916 5302
rect 9770 5264 9826 5273
rect 9864 5238 9916 5244
rect 9770 5199 9826 5208
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9600 4950 9720 4978
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9272 4100 9444 4128
rect 9220 4082 9272 4088
rect 9508 4078 9536 4218
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9600 3890 9628 4950
rect 9678 4856 9734 4865
rect 9734 4814 9812 4842
rect 9876 4826 9904 5034
rect 9678 4791 9734 4800
rect 9678 4720 9734 4729
rect 9678 4655 9734 4664
rect 9692 4146 9720 4655
rect 9784 4554 9812 4814
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9784 4078 9812 4218
rect 9968 4162 9996 5034
rect 9876 4134 9996 4162
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9600 3862 9720 3890
rect 9126 3768 9182 3777
rect 9182 3726 9260 3754
rect 9126 3703 9182 3712
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 9232 3346 9260 3726
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9310 3360 9366 3369
rect 9232 3318 9310 3346
rect 8846 3292 9154 3301
rect 9310 3295 9366 3304
rect 8846 3290 8852 3292
rect 8908 3290 8932 3292
rect 8988 3290 9012 3292
rect 9068 3290 9092 3292
rect 9148 3290 9154 3292
rect 8908 3238 8910 3290
rect 9090 3238 9092 3290
rect 8846 3236 8852 3238
rect 8908 3236 8932 3238
rect 8988 3236 9012 3238
rect 9068 3236 9092 3238
rect 9148 3236 9154 3238
rect 8846 3227 9154 3236
rect 9310 3224 9366 3233
rect 9232 3182 9310 3210
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8758 2408 8814 2417
rect 8576 2032 8628 2038
rect 8576 1974 8628 1980
rect 8576 1828 8628 1834
rect 8576 1770 8628 1776
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 8392 1352 8444 1358
rect 8392 1294 8444 1300
rect 8484 1352 8536 1358
rect 8484 1294 8536 1300
rect 8404 950 8432 1294
rect 8392 944 8444 950
rect 8392 886 8444 892
rect 8496 814 8524 1294
rect 8588 1193 8616 1770
rect 8680 1290 8708 2382
rect 8758 2343 8814 2352
rect 8772 1329 8800 2343
rect 8864 2310 8892 2518
rect 9048 2446 9076 3062
rect 9232 2446 9260 3182
rect 9310 3159 9366 3168
rect 9508 3126 9536 3470
rect 9496 3120 9548 3126
rect 9402 3088 9458 3097
rect 9496 3062 9548 3068
rect 9402 3023 9458 3032
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9324 2666 9352 2926
rect 9416 2774 9444 3023
rect 9692 2922 9720 3862
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9784 3058 9812 3130
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9876 2774 9904 4134
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9968 3194 9996 3606
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10060 3126 10088 5494
rect 10244 5284 10272 5494
rect 10152 5256 10272 5284
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 9416 2746 9536 2774
rect 9324 2638 9444 2666
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9310 2272 9366 2281
rect 8846 2204 9154 2213
rect 8846 2202 8852 2204
rect 8908 2202 8932 2204
rect 8988 2202 9012 2204
rect 9068 2202 9092 2204
rect 9148 2202 9154 2204
rect 8908 2150 8910 2202
rect 9090 2150 9092 2202
rect 8846 2148 8852 2150
rect 8908 2148 8932 2150
rect 8988 2148 9012 2150
rect 9068 2148 9092 2150
rect 9148 2148 9154 2150
rect 8846 2139 9154 2148
rect 9036 2032 9088 2038
rect 9036 1974 9088 1980
rect 8944 1556 8996 1562
rect 8944 1498 8996 1504
rect 8758 1320 8814 1329
rect 8668 1284 8720 1290
rect 8956 1290 8984 1498
rect 9048 1358 9076 1974
rect 9128 1760 9180 1766
rect 9128 1702 9180 1708
rect 9140 1494 9168 1702
rect 9128 1488 9180 1494
rect 9232 1465 9260 2246
rect 9310 2207 9366 2216
rect 9324 1766 9352 2207
rect 9312 1760 9364 1766
rect 9312 1702 9364 1708
rect 9128 1430 9180 1436
rect 9218 1456 9274 1465
rect 9218 1391 9274 1400
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 8758 1255 8814 1264
rect 8944 1284 8996 1290
rect 8668 1226 8720 1232
rect 8944 1226 8996 1232
rect 8574 1184 8630 1193
rect 8574 1119 8630 1128
rect 8846 1116 9154 1125
rect 8846 1114 8852 1116
rect 8908 1114 8932 1116
rect 8988 1114 9012 1116
rect 9068 1114 9092 1116
rect 9148 1114 9154 1116
rect 8908 1062 8910 1114
rect 9090 1062 9092 1114
rect 8846 1060 8852 1062
rect 8908 1060 8932 1062
rect 8988 1060 9012 1062
rect 9068 1060 9092 1062
rect 9148 1060 9154 1062
rect 8846 1051 9154 1060
rect 8484 808 8536 814
rect 7930 776 7986 785
rect 7930 711 7986 720
rect 8206 776 8262 785
rect 8484 750 8536 756
rect 8206 711 8262 720
rect 9416 406 9444 2638
rect 9508 2394 9536 2746
rect 9784 2746 9904 2774
rect 9508 2366 9628 2394
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9508 1562 9536 2246
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 9508 1057 9536 1498
rect 9494 1048 9550 1057
rect 9494 983 9550 992
rect 9600 814 9628 2366
rect 9784 2292 9812 2746
rect 10152 2650 10180 5256
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10244 4729 10272 5102
rect 10336 5098 10364 5902
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 10428 4758 10456 6072
rect 10506 5944 10562 5953
rect 10506 5879 10562 5888
rect 10520 5846 10548 5879
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10506 5672 10562 5681
rect 10506 5607 10562 5616
rect 10520 5352 10548 5607
rect 10612 5545 10640 7262
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10820 7100 11128 7109
rect 10820 7098 10826 7100
rect 10882 7098 10906 7100
rect 10962 7098 10986 7100
rect 11042 7098 11066 7100
rect 11122 7098 11128 7100
rect 10882 7046 10884 7098
rect 11064 7046 11066 7098
rect 10820 7044 10826 7046
rect 10882 7044 10906 7046
rect 10962 7044 10986 7046
rect 11042 7044 11066 7046
rect 11122 7044 11128 7046
rect 10820 7035 11128 7044
rect 11058 6896 11114 6905
rect 11058 6831 11114 6840
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10796 6662 10824 6734
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10784 6656 10836 6662
rect 10888 6633 10916 6734
rect 11072 6633 11100 6831
rect 10784 6598 10836 6604
rect 10874 6624 10930 6633
rect 10598 5536 10654 5545
rect 10598 5471 10654 5480
rect 10520 5324 10640 5352
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10416 4752 10468 4758
rect 10230 4720 10286 4729
rect 10416 4694 10468 4700
rect 10230 4655 10286 4664
rect 10232 4616 10284 4622
rect 10520 4570 10548 5170
rect 10612 5098 10640 5324
rect 10704 5302 10732 6598
rect 10874 6559 10930 6568
rect 11058 6624 11114 6633
rect 11058 6559 11114 6568
rect 11164 6440 11192 8842
rect 11256 8265 11284 9522
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11348 9217 11376 9454
rect 11334 9208 11390 9217
rect 11334 9143 11390 9152
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11348 8786 11376 9046
rect 11440 8906 11468 9862
rect 11624 9674 11652 11614
rect 11702 11520 11758 11529
rect 11702 11455 11758 11464
rect 11532 9646 11652 9674
rect 11532 9450 11560 9646
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11520 9444 11572 9450
rect 11520 9386 11572 9392
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11348 8758 11560 8786
rect 11336 8424 11388 8430
rect 11388 8372 11468 8378
rect 11336 8366 11468 8372
rect 11348 8350 11468 8366
rect 11336 8288 11388 8294
rect 11242 8256 11298 8265
rect 11336 8230 11388 8236
rect 11242 8191 11298 8200
rect 11348 7954 11376 8230
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11440 7857 11468 8350
rect 11532 8294 11560 8758
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11426 7848 11482 7857
rect 11426 7783 11482 7792
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11520 7744 11572 7750
rect 11624 7732 11652 9522
rect 11572 7704 11652 7732
rect 11520 7686 11572 7692
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11256 7041 11284 7278
rect 11242 7032 11298 7041
rect 11242 6967 11298 6976
rect 11072 6412 11192 6440
rect 11072 6361 11100 6412
rect 11058 6352 11114 6361
rect 11058 6287 11114 6296
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 10820 6012 11128 6021
rect 10820 6010 10826 6012
rect 10882 6010 10906 6012
rect 10962 6010 10986 6012
rect 11042 6010 11066 6012
rect 11122 6010 11128 6012
rect 10882 5958 10884 6010
rect 11064 5958 11066 6010
rect 10820 5956 10826 5958
rect 10882 5956 10906 5958
rect 10962 5956 10986 5958
rect 11042 5956 11066 5958
rect 11122 5956 11128 5958
rect 10820 5947 11128 5956
rect 11058 5808 11114 5817
rect 10784 5772 10836 5778
rect 11058 5743 11114 5752
rect 10784 5714 10836 5720
rect 10796 5681 10824 5714
rect 10782 5672 10838 5681
rect 10782 5607 10838 5616
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10796 5166 10824 5306
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10600 5092 10652 5098
rect 10600 5034 10652 5040
rect 11072 5012 11100 5743
rect 11164 5080 11192 6258
rect 11256 5234 11284 6967
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11164 5052 11284 5080
rect 11072 4984 11192 5012
rect 10820 4924 11128 4933
rect 10820 4922 10826 4924
rect 10882 4922 10906 4924
rect 10962 4922 10986 4924
rect 11042 4922 11066 4924
rect 11122 4922 11128 4924
rect 10882 4870 10884 4922
rect 11064 4870 11066 4922
rect 10820 4868 10826 4870
rect 10882 4868 10906 4870
rect 10962 4868 10986 4870
rect 11042 4868 11066 4870
rect 11122 4868 11128 4870
rect 10598 4856 10654 4865
rect 10820 4859 11128 4868
rect 11164 4808 11192 4984
rect 10654 4800 11008 4808
rect 10598 4791 11008 4800
rect 10612 4780 11008 4791
rect 10980 4622 11008 4780
rect 11072 4780 11192 4808
rect 10232 4558 10284 4564
rect 10244 3602 10272 4558
rect 10336 4542 10548 4570
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10230 3224 10286 3233
rect 10230 3159 10286 3168
rect 10244 2825 10272 3159
rect 10230 2816 10286 2825
rect 10230 2751 10286 2760
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 9864 2440 9916 2446
rect 10152 2394 10180 2586
rect 9864 2382 9916 2388
rect 9692 2264 9812 2292
rect 9692 1970 9720 2264
rect 9876 2145 9904 2382
rect 9968 2366 10180 2394
rect 9862 2136 9918 2145
rect 9772 2100 9824 2106
rect 9862 2071 9918 2080
rect 9772 2042 9824 2048
rect 9680 1964 9732 1970
rect 9680 1906 9732 1912
rect 9588 808 9640 814
rect 9588 750 9640 756
rect 9692 678 9720 1906
rect 9784 1902 9812 2042
rect 9876 1970 9904 2071
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 9772 1896 9824 1902
rect 9772 1838 9824 1844
rect 9876 1442 9904 1906
rect 9968 1562 9996 2366
rect 10048 2304 10100 2310
rect 10232 2304 10284 2310
rect 10048 2246 10100 2252
rect 10152 2264 10232 2292
rect 10060 2106 10088 2246
rect 10048 2100 10100 2106
rect 10048 2042 10100 2048
rect 10152 1873 10180 2264
rect 10232 2246 10284 2252
rect 10232 2032 10284 2038
rect 10232 1974 10284 1980
rect 10138 1864 10194 1873
rect 10138 1799 10194 1808
rect 10244 1601 10272 1974
rect 10230 1592 10286 1601
rect 9956 1556 10008 1562
rect 10230 1527 10286 1536
rect 9956 1498 10008 1504
rect 9876 1414 9996 1442
rect 9968 1329 9996 1414
rect 9954 1320 10010 1329
rect 9864 1284 9916 1290
rect 9954 1255 10010 1264
rect 9864 1226 9916 1232
rect 9876 950 9904 1226
rect 10232 1216 10284 1222
rect 10232 1158 10284 1164
rect 9864 944 9916 950
rect 9864 886 9916 892
rect 9680 672 9732 678
rect 9680 614 9732 620
rect 9692 513 9720 614
rect 9678 504 9734 513
rect 9678 439 9734 448
rect 9404 400 9456 406
rect 9404 342 9456 348
rect 9876 270 9904 886
rect 10244 678 10272 1158
rect 10336 746 10364 4542
rect 10690 4312 10746 4321
rect 10690 4247 10746 4256
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10506 3904 10562 3913
rect 10506 3839 10562 3848
rect 10520 3194 10548 3839
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10428 1018 10456 2790
rect 10520 2258 10548 2790
rect 10612 2378 10640 4014
rect 10704 2650 10732 4247
rect 10796 4078 10824 4558
rect 11072 4282 11100 4780
rect 11256 4740 11284 5052
rect 11164 4712 11284 4740
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10980 3924 11008 4218
rect 11164 4078 11192 4712
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11256 4321 11284 4422
rect 11242 4312 11298 4321
rect 11242 4247 11298 4256
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 10980 3896 11192 3924
rect 10820 3836 11128 3845
rect 10820 3834 10826 3836
rect 10882 3834 10906 3836
rect 10962 3834 10986 3836
rect 11042 3834 11066 3836
rect 11122 3834 11128 3836
rect 10882 3782 10884 3834
rect 11064 3782 11066 3834
rect 10820 3780 10826 3782
rect 10882 3780 10906 3782
rect 10962 3780 10986 3782
rect 11042 3780 11066 3782
rect 11122 3780 11128 3782
rect 10820 3771 11128 3780
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10796 2854 10824 3402
rect 10888 3194 10916 3402
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10980 3097 11008 3674
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 10966 3088 11022 3097
rect 10966 3023 11022 3032
rect 10784 2848 10836 2854
rect 10980 2836 11008 3023
rect 11072 2990 11100 3538
rect 11164 3398 11192 3896
rect 11242 3904 11298 3913
rect 11242 3839 11298 3848
rect 11256 3534 11284 3839
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11244 2848 11296 2854
rect 10980 2808 11192 2836
rect 10784 2790 10836 2796
rect 10820 2748 11128 2757
rect 10820 2746 10826 2748
rect 10882 2746 10906 2748
rect 10962 2746 10986 2748
rect 11042 2746 11066 2748
rect 11122 2746 11128 2748
rect 10882 2694 10884 2746
rect 11064 2694 11066 2746
rect 10820 2692 10826 2694
rect 10882 2692 10906 2694
rect 10962 2692 10986 2694
rect 11042 2692 11066 2694
rect 11122 2692 11128 2694
rect 10820 2683 11128 2692
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 11060 2576 11112 2582
rect 10874 2544 10930 2553
rect 11060 2518 11112 2524
rect 10874 2479 10930 2488
rect 10784 2440 10836 2446
rect 10888 2428 10916 2479
rect 10836 2400 10916 2428
rect 10784 2382 10836 2388
rect 10600 2372 10652 2378
rect 10600 2314 10652 2320
rect 11072 2310 11100 2518
rect 10968 2304 11020 2310
rect 10520 2230 10732 2258
rect 10968 2246 11020 2252
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 10704 1902 10732 2230
rect 10782 2136 10838 2145
rect 10782 2071 10838 2080
rect 10796 1970 10824 2071
rect 10876 2032 10928 2038
rect 10876 1974 10928 1980
rect 10784 1964 10836 1970
rect 10784 1906 10836 1912
rect 10692 1896 10744 1902
rect 10888 1873 10916 1974
rect 10692 1838 10744 1844
rect 10874 1864 10930 1873
rect 10508 1828 10560 1834
rect 10508 1770 10560 1776
rect 10520 1562 10548 1770
rect 10508 1556 10560 1562
rect 10508 1498 10560 1504
rect 10508 1284 10560 1290
rect 10508 1226 10560 1232
rect 10520 1018 10548 1226
rect 10416 1012 10468 1018
rect 10416 954 10468 960
rect 10508 1012 10560 1018
rect 10508 954 10560 960
rect 10324 740 10376 746
rect 10324 682 10376 688
rect 10232 672 10284 678
rect 10232 614 10284 620
rect 10704 610 10732 1838
rect 10874 1799 10930 1808
rect 10980 1766 11008 2246
rect 11164 1970 11192 2808
rect 11244 2790 11296 2796
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 10968 1760 11020 1766
rect 10968 1702 11020 1708
rect 10820 1660 11128 1669
rect 10820 1658 10826 1660
rect 10882 1658 10906 1660
rect 10962 1658 10986 1660
rect 11042 1658 11066 1660
rect 11122 1658 11128 1660
rect 10882 1606 10884 1658
rect 11064 1606 11066 1658
rect 10820 1604 10826 1606
rect 10882 1604 10906 1606
rect 10962 1604 10986 1606
rect 11042 1604 11066 1606
rect 11122 1604 11128 1606
rect 10820 1595 11128 1604
rect 11256 1358 11284 2790
rect 11348 2038 11376 7686
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11440 7002 11468 7482
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11440 5574 11468 6666
rect 11532 6390 11560 7686
rect 11610 7304 11666 7313
rect 11610 7239 11612 7248
rect 11664 7239 11666 7248
rect 11612 7210 11664 7216
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11520 6384 11572 6390
rect 11624 6361 11652 6734
rect 11520 6326 11572 6332
rect 11610 6352 11666 6361
rect 11610 6287 11666 6296
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11440 3534 11468 5510
rect 11532 4214 11560 6190
rect 11610 5944 11666 5953
rect 11610 5879 11666 5888
rect 11624 5642 11652 5879
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11610 4992 11666 5001
rect 11610 4927 11666 4936
rect 11624 4214 11652 4927
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11716 3754 11744 11455
rect 11808 10962 11836 12407
rect 11900 11054 11928 14198
rect 11992 11354 12020 15302
rect 12084 15201 12112 18527
rect 12440 18148 12492 18154
rect 12440 18090 12492 18096
rect 12346 17232 12402 17241
rect 12346 17167 12402 17176
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12176 15706 12204 16186
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12162 15328 12218 15337
rect 12162 15263 12218 15272
rect 12070 15192 12126 15201
rect 12070 15127 12126 15136
rect 12070 14920 12126 14929
rect 12070 14855 12126 14864
rect 12084 14618 12112 14855
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12176 14414 12204 15263
rect 12268 15162 12296 15506
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12360 15008 12388 17167
rect 12452 15026 12480 18090
rect 12544 15638 12572 19790
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 12794 19612 13102 19621
rect 12794 19610 12800 19612
rect 12856 19610 12880 19612
rect 12936 19610 12960 19612
rect 13016 19610 13040 19612
rect 13096 19610 13102 19612
rect 12856 19558 12858 19610
rect 13038 19558 13040 19610
rect 12794 19556 12800 19558
rect 12856 19556 12880 19558
rect 12936 19556 12960 19558
rect 13016 19556 13040 19558
rect 13096 19556 13102 19558
rect 12794 19547 13102 19556
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 12794 18524 13102 18533
rect 12794 18522 12800 18524
rect 12856 18522 12880 18524
rect 12936 18522 12960 18524
rect 13016 18522 13040 18524
rect 13096 18522 13102 18524
rect 12856 18470 12858 18522
rect 13038 18470 13040 18522
rect 12794 18468 12800 18470
rect 12856 18468 12880 18470
rect 12936 18468 12960 18470
rect 13016 18468 13040 18470
rect 13096 18468 13102 18470
rect 12794 18459 13102 18468
rect 12794 17436 13102 17445
rect 12794 17434 12800 17436
rect 12856 17434 12880 17436
rect 12936 17434 12960 17436
rect 13016 17434 13040 17436
rect 13096 17434 13102 17436
rect 12856 17382 12858 17434
rect 13038 17382 13040 17434
rect 12794 17380 12800 17382
rect 12856 17380 12880 17382
rect 12936 17380 12960 17382
rect 13016 17380 13040 17382
rect 13096 17380 13102 17382
rect 12794 17371 13102 17380
rect 12794 16348 13102 16357
rect 12794 16346 12800 16348
rect 12856 16346 12880 16348
rect 12936 16346 12960 16348
rect 13016 16346 13040 16348
rect 13096 16346 13102 16348
rect 12856 16294 12858 16346
rect 13038 16294 13040 16346
rect 12794 16292 12800 16294
rect 12856 16292 12880 16294
rect 12936 16292 12960 16294
rect 13016 16292 13040 16294
rect 13096 16292 13102 16294
rect 12794 16283 13102 16292
rect 13082 16144 13138 16153
rect 13082 16079 13138 16088
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12532 15632 12584 15638
rect 12532 15574 12584 15580
rect 12268 14980 12388 15008
rect 12440 15020 12492 15026
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12162 14240 12218 14249
rect 12162 14175 12218 14184
rect 12070 14104 12126 14113
rect 12070 14039 12126 14048
rect 12084 14006 12112 14039
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12084 13705 12112 13806
rect 12070 13696 12126 13705
rect 12070 13631 12126 13640
rect 12176 13530 12204 14175
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 12162 13288 12218 13297
rect 12162 13223 12218 13232
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12084 12764 12112 13126
rect 12176 12832 12204 13223
rect 12268 12986 12296 14980
rect 12440 14962 12492 14968
rect 12544 14906 12572 15574
rect 12636 14929 12664 15914
rect 13096 15706 13124 16079
rect 13174 15872 13230 15881
rect 13174 15807 13230 15816
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 12898 15600 12954 15609
rect 12898 15535 12900 15544
rect 12952 15535 12954 15544
rect 12900 15506 12952 15512
rect 12992 15496 13044 15502
rect 12714 15464 12770 15473
rect 12714 15399 12770 15408
rect 12990 15464 12992 15473
rect 13044 15464 13046 15473
rect 12990 15399 13046 15408
rect 12360 14878 12572 14906
rect 12622 14920 12678 14929
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12176 12804 12296 12832
rect 12084 12736 12204 12764
rect 12070 11792 12126 11801
rect 12070 11727 12072 11736
rect 12124 11727 12126 11736
rect 12072 11698 12124 11704
rect 12176 11642 12204 12736
rect 12268 12481 12296 12804
rect 12254 12472 12310 12481
rect 12254 12407 12310 12416
rect 12254 12064 12310 12073
rect 12254 11999 12310 12008
rect 12084 11614 12204 11642
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12084 11150 12112 11614
rect 12268 11540 12296 11999
rect 12360 11937 12388 14878
rect 12622 14855 12678 14864
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12452 13394 12480 14758
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12544 13462 12572 14418
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12532 13320 12584 13326
rect 12530 13288 12532 13297
rect 12584 13288 12586 13297
rect 12530 13223 12586 13232
rect 12438 13152 12494 13161
rect 12494 13110 12572 13138
rect 12438 13087 12494 13096
rect 12438 13016 12494 13025
rect 12438 12951 12494 12960
rect 12452 12753 12480 12951
rect 12544 12850 12572 13110
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12438 12744 12494 12753
rect 12438 12679 12494 12688
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12346 11928 12402 11937
rect 12346 11863 12402 11872
rect 12176 11512 12388 11540
rect 12176 11354 12204 11512
rect 12254 11384 12310 11393
rect 12164 11348 12216 11354
rect 12254 11319 12310 11328
rect 12164 11290 12216 11296
rect 12072 11144 12124 11150
rect 12164 11144 12216 11150
rect 12072 11086 12124 11092
rect 12162 11112 12164 11121
rect 12268 11132 12296 11319
rect 12360 11200 12388 11512
rect 12452 11506 12480 12582
rect 12544 11608 12572 12650
rect 12636 11744 12664 14855
rect 12728 14770 12756 15399
rect 12794 15260 13102 15269
rect 12794 15258 12800 15260
rect 12856 15258 12880 15260
rect 12936 15258 12960 15260
rect 13016 15258 13040 15260
rect 13096 15258 13102 15260
rect 12856 15206 12858 15258
rect 13038 15206 13040 15258
rect 12794 15204 12800 15206
rect 12856 15204 12880 15206
rect 12936 15204 12960 15206
rect 13016 15204 13040 15206
rect 13096 15204 13102 15206
rect 12794 15195 13102 15204
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12728 14742 12848 14770
rect 12714 14648 12770 14657
rect 12714 14583 12770 14592
rect 12728 14482 12756 14583
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12820 14260 12848 14742
rect 12912 14618 12940 14962
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 13188 14414 13216 15807
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 12728 14232 12848 14260
rect 12728 14056 12756 14232
rect 12794 14172 13102 14181
rect 12794 14170 12800 14172
rect 12856 14170 12880 14172
rect 12936 14170 12960 14172
rect 13016 14170 13040 14172
rect 13096 14170 13102 14172
rect 12856 14118 12858 14170
rect 13038 14118 13040 14170
rect 12794 14116 12800 14118
rect 12856 14116 12880 14118
rect 12936 14116 12960 14118
rect 13016 14116 13040 14118
rect 13096 14116 13102 14118
rect 12794 14107 13102 14116
rect 12728 14028 12940 14056
rect 12912 13938 12940 14028
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12728 13841 12756 13874
rect 12808 13864 12860 13870
rect 12714 13832 12770 13841
rect 12808 13806 12860 13812
rect 12714 13767 12770 13776
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12728 11880 12756 13398
rect 12820 13258 12848 13806
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 13530 12940 13670
rect 12990 13560 13046 13569
rect 12900 13524 12952 13530
rect 12990 13495 13046 13504
rect 13096 13512 13124 13874
rect 13176 13524 13228 13530
rect 12900 13466 12952 13472
rect 13004 13394 13032 13495
rect 13096 13484 13176 13512
rect 13176 13466 13228 13472
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12794 13084 13102 13093
rect 12794 13082 12800 13084
rect 12856 13082 12880 13084
rect 12936 13082 12960 13084
rect 13016 13082 13040 13084
rect 13096 13082 13102 13084
rect 12856 13030 12858 13082
rect 13038 13030 13040 13082
rect 12794 13028 12800 13030
rect 12856 13028 12880 13030
rect 12936 13028 12960 13030
rect 13016 13028 13040 13030
rect 13096 13028 13102 13030
rect 12794 13019 13102 13028
rect 12808 12980 12860 12986
rect 13188 12968 13216 13466
rect 12808 12922 12860 12928
rect 13096 12940 13216 12968
rect 12820 12850 12848 12922
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12898 12744 12954 12753
rect 13004 12714 13032 12854
rect 12898 12679 12954 12688
rect 12992 12708 13044 12714
rect 12912 12102 12940 12679
rect 12992 12650 13044 12656
rect 13096 12374 13124 12940
rect 13174 12472 13230 12481
rect 13174 12407 13176 12416
rect 13228 12407 13230 12416
rect 13176 12378 13228 12384
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 13280 12186 13308 14758
rect 13372 12646 13400 15370
rect 13464 14634 13492 18838
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13556 14793 13584 15098
rect 13542 14784 13598 14793
rect 13542 14719 13598 14728
rect 13464 14606 13584 14634
rect 13556 14521 13584 14606
rect 13542 14512 13598 14521
rect 13542 14447 13544 14456
rect 13596 14447 13598 14456
rect 13544 14418 13596 14424
rect 13452 14408 13504 14414
rect 13556 14387 13584 14418
rect 13648 14414 13676 17274
rect 13726 15600 13782 15609
rect 13726 15535 13782 15544
rect 13740 15162 13768 15535
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13832 15026 13860 18770
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13636 14408 13688 14414
rect 13452 14350 13504 14356
rect 13636 14350 13688 14356
rect 13464 14249 13492 14350
rect 13636 14272 13688 14278
rect 13450 14240 13506 14249
rect 13636 14214 13688 14220
rect 13450 14175 13506 14184
rect 13450 13832 13506 13841
rect 13450 13767 13506 13776
rect 13464 13326 13492 13767
rect 13542 13560 13598 13569
rect 13542 13495 13598 13504
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13556 13258 13584 13495
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13450 13016 13506 13025
rect 13450 12951 13506 12960
rect 13464 12918 13492 12951
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13648 12434 13676 14214
rect 13740 13569 13768 14962
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13726 13560 13782 13569
rect 13726 13495 13782 13504
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13188 12158 13308 12186
rect 13372 12406 13676 12434
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12794 11996 13102 12005
rect 12794 11994 12800 11996
rect 12856 11994 12880 11996
rect 12936 11994 12960 11996
rect 13016 11994 13040 11996
rect 13096 11994 13102 11996
rect 12856 11942 12858 11994
rect 13038 11942 13040 11994
rect 12794 11940 12800 11942
rect 12856 11940 12880 11942
rect 12936 11940 12960 11942
rect 13016 11940 13040 11942
rect 13096 11940 13102 11942
rect 12794 11931 13102 11940
rect 12728 11852 12940 11880
rect 12716 11756 12768 11762
rect 12636 11716 12716 11744
rect 12716 11698 12768 11704
rect 12544 11580 12848 11608
rect 12452 11478 12756 11506
rect 12530 11384 12586 11393
rect 12530 11319 12586 11328
rect 12624 11348 12676 11354
rect 12360 11172 12480 11200
rect 12216 11112 12218 11121
rect 12268 11104 12388 11132
rect 11900 11026 12112 11054
rect 12162 11047 12218 11056
rect 12084 10996 12112 11026
rect 12084 10968 12204 10996
rect 11808 10934 11928 10962
rect 11794 9616 11850 9625
rect 11794 9551 11850 9560
rect 11808 4214 11836 9551
rect 11900 7857 11928 10934
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11992 9761 12020 10202
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 11978 9752 12034 9761
rect 11978 9687 12034 9696
rect 11980 9648 12032 9654
rect 11978 9616 11980 9625
rect 12032 9616 12034 9625
rect 11978 9551 12034 9560
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11992 8090 12020 8842
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11886 7848 11942 7857
rect 11886 7783 11942 7792
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11992 7478 12020 7686
rect 12084 7546 12112 9998
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 11980 7472 12032 7478
rect 12176 7426 12204 10968
rect 12254 10840 12310 10849
rect 12254 10775 12310 10784
rect 12268 10470 12296 10775
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12360 10282 12388 11104
rect 12452 10470 12480 11172
rect 12544 10810 12572 11319
rect 12624 11290 12676 11296
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 11980 7414 12032 7420
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 12084 7398 12204 7426
rect 12268 10254 12388 10282
rect 11900 5914 11928 7346
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11992 6662 12020 7278
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11978 6488 12034 6497
rect 11978 6423 12034 6432
rect 11992 6390 12020 6423
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11886 5808 11942 5817
rect 11886 5743 11888 5752
rect 11940 5743 11942 5752
rect 11888 5714 11940 5720
rect 12084 5574 12112 7398
rect 12268 6798 12296 10254
rect 12544 10062 12572 10542
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12530 9888 12586 9897
rect 12530 9823 12586 9832
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12360 9353 12388 9522
rect 12544 9450 12572 9823
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12346 9344 12402 9353
rect 12346 9279 12402 9288
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12544 8945 12572 9046
rect 12530 8936 12586 8945
rect 12348 8900 12400 8906
rect 12530 8871 12586 8880
rect 12348 8842 12400 8848
rect 12360 8498 12388 8842
rect 12530 8664 12586 8673
rect 12440 8628 12492 8634
rect 12530 8599 12586 8608
rect 12440 8570 12492 8576
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12360 6644 12388 7890
rect 12452 7857 12480 8570
rect 12438 7848 12494 7857
rect 12438 7783 12494 7792
rect 12438 7712 12494 7721
rect 12438 7647 12494 7656
rect 12452 7290 12480 7647
rect 12544 7478 12572 8599
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12452 7262 12572 7290
rect 12438 7168 12494 7177
rect 12438 7103 12494 7112
rect 12268 6616 12388 6644
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12072 5568 12124 5574
rect 11886 5536 11942 5545
rect 11942 5494 12020 5522
rect 12072 5510 12124 5516
rect 11886 5471 11942 5480
rect 11886 5400 11942 5409
rect 11886 5335 11942 5344
rect 11900 5098 11928 5335
rect 11992 5234 12020 5494
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 12084 4826 12112 5510
rect 12176 5409 12204 6054
rect 12162 5400 12218 5409
rect 12162 5335 12218 5344
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12176 5137 12204 5170
rect 12162 5128 12218 5137
rect 12162 5063 12218 5072
rect 12268 5030 12296 6616
rect 12452 6372 12480 7103
rect 12544 6866 12572 7262
rect 12636 6934 12664 11290
rect 12728 9704 12756 11478
rect 12820 11354 12848 11580
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12912 11234 12940 11852
rect 13188 11830 13216 12158
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11898 13308 12038
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13268 11620 13320 11626
rect 12820 11206 12940 11234
rect 13004 11580 13268 11608
rect 12820 11150 12848 11206
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 13004 11014 13032 11580
rect 13268 11562 13320 11568
rect 13372 11370 13400 12406
rect 13452 12368 13504 12374
rect 13450 12336 13452 12345
rect 13504 12336 13506 12345
rect 13740 12322 13768 13126
rect 13832 12889 13860 14214
rect 13924 14006 13952 18906
rect 14016 14414 14044 19654
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 14002 14104 14058 14113
rect 14002 14039 14004 14048
rect 14056 14039 14058 14048
rect 14004 14010 14056 14016
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 14002 13968 14058 13977
rect 14002 13903 14058 13912
rect 14016 13870 14044 13903
rect 14004 13864 14056 13870
rect 13910 13832 13966 13841
rect 14004 13806 14056 13812
rect 13910 13767 13966 13776
rect 13818 12880 13874 12889
rect 13818 12815 13874 12824
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13450 12271 13506 12280
rect 13556 12294 13768 12322
rect 13450 11928 13506 11937
rect 13450 11863 13506 11872
rect 13464 11830 13492 11863
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13556 11642 13584 12294
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13648 11880 13676 12174
rect 13726 12064 13782 12073
rect 13726 11999 13782 12008
rect 13740 11898 13768 11999
rect 13832 11914 13860 12582
rect 13924 12306 13952 13767
rect 14002 13696 14058 13705
rect 14002 13631 14058 13640
rect 14016 12918 14044 13631
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 14108 12850 14136 16118
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14200 13705 14228 14894
rect 14292 14618 14320 16934
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14186 13696 14242 13705
rect 14186 13631 14242 13640
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14200 13025 14228 13126
rect 14186 13016 14242 13025
rect 14186 12951 14242 12960
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14186 12744 14242 12753
rect 14004 12708 14056 12714
rect 14186 12679 14242 12688
rect 14004 12650 14056 12656
rect 14016 12617 14044 12650
rect 14096 12640 14148 12646
rect 14002 12608 14058 12617
rect 14148 12588 14156 12594
rect 14096 12582 14156 12588
rect 14108 12566 14156 12582
rect 14002 12543 14058 12552
rect 14128 12442 14156 12566
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14096 12436 14156 12442
rect 14148 12396 14156 12436
rect 14096 12378 14148 12384
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13645 11852 13676 11880
rect 13728 11892 13780 11898
rect 13645 11778 13673 11852
rect 13832 11886 13952 11914
rect 13728 11834 13780 11840
rect 13924 11812 13952 11886
rect 14016 11880 14044 12378
rect 14094 12336 14150 12345
rect 14094 12271 14096 12280
rect 14148 12271 14150 12280
rect 14096 12242 14148 12248
rect 14016 11852 14136 11880
rect 13924 11784 14044 11812
rect 13645 11750 13676 11778
rect 13648 11744 13676 11750
rect 13648 11716 13952 11744
rect 13556 11614 13768 11642
rect 13740 11529 13768 11614
rect 13820 11552 13872 11558
rect 13726 11520 13782 11529
rect 13820 11494 13872 11500
rect 13726 11455 13782 11464
rect 13096 11342 13400 11370
rect 13096 11150 13124 11342
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12794 10908 13102 10917
rect 12794 10906 12800 10908
rect 12856 10906 12880 10908
rect 12936 10906 12960 10908
rect 13016 10906 13040 10908
rect 13096 10906 13102 10908
rect 12856 10854 12858 10906
rect 13038 10854 13040 10906
rect 12794 10852 12800 10854
rect 12856 10852 12880 10854
rect 12936 10852 12960 10854
rect 13016 10852 13040 10854
rect 13096 10852 13102 10854
rect 12794 10843 13102 10852
rect 13188 10810 13216 11222
rect 13372 11098 13400 11342
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13372 11070 13492 11098
rect 13360 11008 13412 11014
rect 13266 10976 13322 10985
rect 13360 10950 13412 10956
rect 13464 10962 13492 11070
rect 13648 11054 13676 11154
rect 13740 11150 13768 11455
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13628 11026 13676 11054
rect 13628 10962 13656 11026
rect 13266 10911 13322 10920
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12820 10577 12848 10610
rect 12806 10568 12862 10577
rect 12806 10503 12862 10512
rect 13174 10568 13230 10577
rect 13174 10503 13230 10512
rect 12820 10266 12848 10503
rect 13188 10470 13216 10503
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13280 10282 13308 10911
rect 13372 10441 13400 10950
rect 13464 10934 13656 10962
rect 13832 10826 13860 11494
rect 13648 10798 13860 10826
rect 13648 10792 13676 10798
rect 13556 10764 13676 10792
rect 13556 10554 13584 10764
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13464 10538 13584 10554
rect 13452 10532 13584 10538
rect 13504 10526 13584 10532
rect 13452 10474 13504 10480
rect 13544 10464 13596 10470
rect 13358 10432 13414 10441
rect 13544 10406 13596 10412
rect 13358 10367 13414 10376
rect 13450 10296 13506 10305
rect 12808 10260 12860 10266
rect 13280 10254 13400 10282
rect 12808 10202 12860 10208
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 12808 10056 12860 10062
rect 12992 10056 13044 10062
rect 12808 9998 12860 10004
rect 12990 10024 12992 10033
rect 13044 10024 13046 10033
rect 12820 9908 12848 9998
rect 12990 9959 13046 9968
rect 12820 9880 13216 9908
rect 12794 9820 13102 9829
rect 12794 9818 12800 9820
rect 12856 9818 12880 9820
rect 12936 9818 12960 9820
rect 13016 9818 13040 9820
rect 13096 9818 13102 9820
rect 12856 9766 12858 9818
rect 13038 9766 13040 9818
rect 12794 9764 12800 9766
rect 12856 9764 12880 9766
rect 12936 9764 12960 9766
rect 13016 9764 13040 9766
rect 13096 9764 13102 9766
rect 12794 9755 13102 9764
rect 13188 9704 13216 9880
rect 13280 9722 13308 10066
rect 12728 9676 12848 9704
rect 12820 9110 12848 9676
rect 13096 9676 13216 9704
rect 13268 9716 13320 9722
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12912 9450 12940 9590
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12728 7993 12756 8978
rect 12992 8968 13044 8974
rect 12990 8936 12992 8945
rect 13044 8936 13046 8945
rect 12990 8871 13046 8880
rect 13096 8820 13124 9676
rect 13268 9658 13320 9664
rect 13372 9602 13400 10254
rect 13450 10231 13506 10240
rect 13464 9897 13492 10231
rect 13450 9888 13506 9897
rect 13450 9823 13506 9832
rect 13372 9574 13492 9602
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13266 9072 13322 9081
rect 13266 9007 13322 9016
rect 13096 8792 13216 8820
rect 12794 8732 13102 8741
rect 12794 8730 12800 8732
rect 12856 8730 12880 8732
rect 12936 8730 12960 8732
rect 13016 8730 13040 8732
rect 13096 8730 13102 8732
rect 12856 8678 12858 8730
rect 13038 8678 13040 8730
rect 12794 8676 12800 8678
rect 12856 8676 12880 8678
rect 12936 8676 12960 8678
rect 13016 8676 13040 8678
rect 13096 8676 13102 8678
rect 12794 8667 13102 8676
rect 13188 8616 13216 8792
rect 13096 8588 13216 8616
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12714 7984 12770 7993
rect 12714 7919 12770 7928
rect 12820 7732 12848 8434
rect 12912 7993 12940 8502
rect 13096 8362 13124 8588
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 12898 7984 12954 7993
rect 12898 7919 12954 7928
rect 12728 7704 12848 7732
rect 12728 7206 12756 7704
rect 12794 7644 13102 7653
rect 12794 7642 12800 7644
rect 12856 7642 12880 7644
rect 12936 7642 12960 7644
rect 13016 7642 13040 7644
rect 13096 7642 13102 7644
rect 12856 7590 12858 7642
rect 13038 7590 13040 7642
rect 12794 7588 12800 7590
rect 12856 7588 12880 7590
rect 12936 7588 12960 7590
rect 13016 7588 13040 7590
rect 13096 7588 13102 7590
rect 12794 7579 13102 7588
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12820 6746 12848 7210
rect 12912 6798 12940 7482
rect 13280 7460 13308 9007
rect 13372 8022 13400 9454
rect 13464 8634 13492 9574
rect 13556 8634 13584 10406
rect 13648 9994 13676 10610
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13634 9480 13690 9489
rect 13634 9415 13690 9424
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13648 8480 13676 9415
rect 13740 8974 13768 10678
rect 13924 10441 13952 11716
rect 14016 10985 14044 11784
rect 14108 11694 14136 11852
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 14200 11558 14228 12679
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14108 11234 14136 11290
rect 14108 11206 14156 11234
rect 14128 11150 14156 11206
rect 14096 11144 14156 11150
rect 14148 11104 14156 11144
rect 14096 11086 14148 11092
rect 14002 10976 14058 10985
rect 14002 10911 14058 10920
rect 14108 10792 14136 11086
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14200 10810 14228 10950
rect 14016 10764 14136 10792
rect 14188 10804 14240 10810
rect 13910 10432 13966 10441
rect 13910 10367 13966 10376
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13740 8673 13768 8910
rect 13726 8664 13782 8673
rect 13726 8599 13782 8608
rect 13728 8560 13780 8566
rect 13464 8452 13676 8480
rect 13726 8528 13728 8537
rect 13780 8528 13782 8537
rect 13726 8463 13782 8472
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13464 7886 13492 8452
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13556 8022 13584 8298
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13360 7472 13412 7478
rect 13280 7432 13360 7460
rect 13360 7414 13412 7420
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12544 6718 12848 6746
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12544 6662 12572 6718
rect 12532 6656 12584 6662
rect 13004 6644 13032 7346
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 12636 6633 13032 6644
rect 12532 6598 12584 6604
rect 12622 6624 13032 6633
rect 12678 6616 13032 6624
rect 12622 6559 12678 6568
rect 12794 6556 13102 6565
rect 12794 6554 12800 6556
rect 12856 6554 12880 6556
rect 12936 6554 12960 6556
rect 13016 6554 13040 6556
rect 13096 6554 13102 6556
rect 12856 6502 12858 6554
rect 13038 6502 13040 6554
rect 12794 6500 12800 6502
rect 12856 6500 12880 6502
rect 12936 6500 12960 6502
rect 13016 6500 13040 6502
rect 13096 6500 13102 6502
rect 12794 6491 13102 6500
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12452 6344 12572 6372
rect 12544 6118 12572 6344
rect 12806 6352 12862 6361
rect 12806 6287 12862 6296
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12360 5234 12388 5850
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12452 5574 12480 5782
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12544 5409 12572 5782
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12530 5400 12586 5409
rect 12530 5335 12586 5344
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12346 5128 12402 5137
rect 12346 5063 12348 5072
rect 12400 5063 12402 5072
rect 12348 5034 12400 5040
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12452 4842 12480 5170
rect 12072 4820 12124 4826
rect 12268 4814 12480 4842
rect 12544 4842 12572 5238
rect 12636 5001 12664 5714
rect 12622 4992 12678 5001
rect 12622 4927 12678 4936
rect 12544 4814 12664 4842
rect 12268 4808 12296 4814
rect 12072 4762 12124 4768
rect 12176 4780 12296 4808
rect 11978 4584 12034 4593
rect 11978 4519 12034 4528
rect 11886 4312 11942 4321
rect 11886 4247 11942 4256
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11624 3726 11744 3754
rect 11900 3738 11928 4247
rect 11888 3732 11940 3738
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11532 3126 11560 3402
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 11624 2774 11652 3726
rect 11888 3674 11940 3680
rect 11704 3664 11756 3670
rect 11702 3632 11704 3641
rect 11756 3632 11758 3641
rect 11702 3567 11758 3576
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 3369 11928 3470
rect 11992 3466 12020 4519
rect 12070 4448 12126 4457
rect 12176 4434 12204 4780
rect 12348 4752 12400 4758
rect 12400 4712 12480 4740
rect 12348 4694 12400 4700
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12126 4406 12204 4434
rect 12070 4383 12126 4392
rect 12268 4214 12296 4490
rect 12452 4282 12480 4712
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12346 4176 12402 4185
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11886 3360 11942 3369
rect 11886 3295 11942 3304
rect 12084 3346 12112 4082
rect 12176 4078 12204 4150
rect 12346 4111 12348 4120
rect 12400 4111 12402 4120
rect 12348 4082 12400 4088
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12256 3936 12308 3942
rect 12308 3896 12388 3924
rect 12256 3878 12308 3884
rect 12360 3738 12388 3896
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 12176 3534 12204 3606
rect 12268 3534 12296 3674
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12256 3528 12308 3534
rect 12308 3488 12388 3516
rect 12256 3470 12308 3476
rect 12084 3318 12296 3346
rect 11702 3088 11758 3097
rect 11702 3023 11758 3032
rect 11440 2746 11652 2774
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11336 1896 11388 1902
rect 11336 1838 11388 1844
rect 11348 1737 11376 1838
rect 11334 1728 11390 1737
rect 11334 1663 11390 1672
rect 11244 1352 11296 1358
rect 11244 1294 11296 1300
rect 11336 1352 11388 1358
rect 11336 1294 11388 1300
rect 10692 604 10744 610
rect 10692 546 10744 552
rect 11348 474 11376 1294
rect 11440 1290 11468 2746
rect 11716 2530 11744 3023
rect 11900 2854 11928 3295
rect 12084 3194 12112 3318
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 12176 2774 12204 3130
rect 11992 2746 12204 2774
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11532 2502 11744 2530
rect 11532 1562 11560 2502
rect 11612 2440 11664 2446
rect 11796 2440 11848 2446
rect 11612 2382 11664 2388
rect 11716 2400 11796 2428
rect 11520 1556 11572 1562
rect 11520 1498 11572 1504
rect 11624 1358 11652 2382
rect 11716 1748 11744 2400
rect 11796 2382 11848 2388
rect 11900 2106 11928 2586
rect 11992 2582 12020 2746
rect 12070 2680 12126 2689
rect 12070 2615 12126 2624
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 12084 2514 12112 2615
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12176 2417 12204 2450
rect 12162 2408 12218 2417
rect 12162 2343 12218 2352
rect 12268 2258 12296 3318
rect 12360 2854 12388 3488
rect 12452 3126 12480 4218
rect 12544 3194 12572 4626
rect 12636 4321 12664 4814
rect 12622 4312 12678 4321
rect 12622 4247 12678 4256
rect 12622 3904 12678 3913
rect 12622 3839 12678 3848
rect 12636 3233 12664 3839
rect 12728 3534 12756 6122
rect 12820 5642 12848 6287
rect 13096 5778 13124 6394
rect 13188 5817 13216 7142
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13280 6633 13308 6938
rect 13464 6905 13492 7822
rect 13450 6896 13506 6905
rect 13450 6831 13506 6840
rect 13360 6792 13412 6798
rect 13556 6780 13584 7958
rect 13412 6752 13584 6780
rect 13360 6734 13412 6740
rect 13266 6624 13322 6633
rect 13266 6559 13322 6568
rect 13372 6322 13400 6734
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13174 5808 13230 5817
rect 13084 5772 13136 5778
rect 13174 5743 13230 5752
rect 13084 5714 13136 5720
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12794 5468 13102 5477
rect 12794 5466 12800 5468
rect 12856 5466 12880 5468
rect 12936 5466 12960 5468
rect 13016 5466 13040 5468
rect 13096 5466 13102 5468
rect 12856 5414 12858 5466
rect 13038 5414 13040 5466
rect 12794 5412 12800 5414
rect 12856 5412 12880 5414
rect 12936 5412 12960 5414
rect 13016 5412 13040 5414
rect 13096 5412 13102 5414
rect 12794 5403 13102 5412
rect 13188 5302 13216 5743
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12820 4865 12848 5034
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 12806 4856 12862 4865
rect 12806 4791 12862 4800
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12820 4622 12848 4694
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12912 4554 12940 4966
rect 13004 4826 13032 4966
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 13280 4740 13308 6054
rect 13372 5817 13400 6258
rect 13464 5914 13492 6598
rect 13542 6488 13598 6497
rect 13542 6423 13598 6432
rect 13556 6118 13584 6423
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13358 5808 13414 5817
rect 13358 5743 13414 5752
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13372 5234 13400 5510
rect 13452 5296 13504 5302
rect 13452 5238 13504 5244
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13188 4712 13308 4740
rect 12900 4548 12952 4554
rect 12900 4490 12952 4496
rect 12794 4380 13102 4389
rect 12794 4378 12800 4380
rect 12856 4378 12880 4380
rect 12936 4378 12960 4380
rect 13016 4378 13040 4380
rect 13096 4378 13102 4380
rect 12856 4326 12858 4378
rect 13038 4326 13040 4378
rect 12794 4324 12800 4326
rect 12856 4324 12880 4326
rect 12936 4324 12960 4326
rect 13016 4324 13040 4326
rect 13096 4324 13102 4326
rect 12794 4315 13102 4324
rect 13188 3913 13216 4712
rect 13360 4616 13412 4622
rect 13280 4576 13360 4604
rect 13280 4214 13308 4576
rect 13360 4558 13412 4564
rect 13464 4486 13492 5238
rect 13556 4593 13584 5714
rect 13542 4584 13598 4593
rect 13542 4519 13598 4528
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13648 4264 13676 8298
rect 13832 7936 13860 9930
rect 13924 8129 13952 10202
rect 14016 9081 14044 10764
rect 14188 10746 14240 10752
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14108 10470 14136 10610
rect 14292 10554 14320 13738
rect 14384 13025 14412 22066
rect 14768 21244 15076 21253
rect 14768 21242 14774 21244
rect 14830 21242 14854 21244
rect 14910 21242 14934 21244
rect 14990 21242 15014 21244
rect 15070 21242 15076 21244
rect 14830 21190 14832 21242
rect 15012 21190 15014 21242
rect 14768 21188 14774 21190
rect 14830 21188 14854 21190
rect 14910 21188 14934 21190
rect 14990 21188 15014 21190
rect 15070 21188 15076 21190
rect 14768 21179 15076 21188
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 14768 20156 15076 20165
rect 14768 20154 14774 20156
rect 14830 20154 14854 20156
rect 14910 20154 14934 20156
rect 14990 20154 15014 20156
rect 15070 20154 15076 20156
rect 14830 20102 14832 20154
rect 15012 20102 15014 20154
rect 14768 20100 14774 20102
rect 14830 20100 14854 20102
rect 14910 20100 14934 20102
rect 14990 20100 15014 20102
rect 15070 20100 15076 20102
rect 14768 20091 15076 20100
rect 14768 19068 15076 19077
rect 14768 19066 14774 19068
rect 14830 19066 14854 19068
rect 14910 19066 14934 19068
rect 14990 19066 15014 19068
rect 15070 19066 15076 19068
rect 14830 19014 14832 19066
rect 15012 19014 15014 19066
rect 14768 19012 14774 19014
rect 14830 19012 14854 19014
rect 14910 19012 14934 19014
rect 14990 19012 15014 19014
rect 15070 19012 15076 19014
rect 14768 19003 15076 19012
rect 15198 18728 15254 18737
rect 15198 18663 15254 18672
rect 14768 17980 15076 17989
rect 14768 17978 14774 17980
rect 14830 17978 14854 17980
rect 14910 17978 14934 17980
rect 14990 17978 15014 17980
rect 15070 17978 15076 17980
rect 14830 17926 14832 17978
rect 15012 17926 15014 17978
rect 14768 17924 14774 17926
rect 14830 17924 14854 17926
rect 14910 17924 14934 17926
rect 14990 17924 15014 17926
rect 15070 17924 15076 17926
rect 14768 17915 15076 17924
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14476 14090 14504 17478
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 14768 16892 15076 16901
rect 14768 16890 14774 16892
rect 14830 16890 14854 16892
rect 14910 16890 14934 16892
rect 14990 16890 15014 16892
rect 15070 16890 15076 16892
rect 14830 16838 14832 16890
rect 15012 16838 15014 16890
rect 14768 16836 14774 16838
rect 14830 16836 14854 16838
rect 14910 16836 14934 16838
rect 14990 16836 15014 16838
rect 15070 16836 15076 16838
rect 14768 16827 15076 16836
rect 14556 16516 14608 16522
rect 14556 16458 14608 16464
rect 14568 15706 14596 16458
rect 14768 15804 15076 15813
rect 14768 15802 14774 15804
rect 14830 15802 14854 15804
rect 14910 15802 14934 15804
rect 14990 15802 15014 15804
rect 15070 15802 15076 15804
rect 14830 15750 14832 15802
rect 15012 15750 15014 15802
rect 14768 15748 14774 15750
rect 14830 15748 14854 15750
rect 14910 15748 14934 15750
rect 14990 15748 15014 15750
rect 15070 15748 15076 15750
rect 14768 15739 15076 15748
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14768 14716 15076 14725
rect 14768 14714 14774 14716
rect 14830 14714 14854 14716
rect 14910 14714 14934 14716
rect 14990 14714 15014 14716
rect 15070 14714 15076 14716
rect 14830 14662 14832 14714
rect 15012 14662 15014 14714
rect 14768 14660 14774 14662
rect 14830 14660 14854 14662
rect 14910 14660 14934 14662
rect 14990 14660 15014 14662
rect 15070 14660 15076 14662
rect 14768 14651 15076 14660
rect 14924 14408 14976 14414
rect 14922 14376 14924 14385
rect 14976 14376 14978 14385
rect 14648 14340 14700 14346
rect 14922 14311 14978 14320
rect 14648 14282 14700 14288
rect 14476 14062 14596 14090
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14476 13705 14504 13942
rect 14568 13841 14596 14062
rect 14554 13832 14610 13841
rect 14554 13767 14610 13776
rect 14462 13696 14518 13705
rect 14462 13631 14518 13640
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14568 13326 14596 13466
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14370 13016 14426 13025
rect 14370 12951 14426 12960
rect 14370 12880 14426 12889
rect 14370 12815 14426 12824
rect 14384 12306 14412 12815
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14370 12200 14426 12209
rect 14370 12135 14426 12144
rect 14384 11830 14412 12135
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14292 10526 14412 10554
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14278 10432 14334 10441
rect 14096 10192 14148 10198
rect 14200 10169 14228 10406
rect 14278 10367 14334 10376
rect 14096 10134 14148 10140
rect 14186 10160 14242 10169
rect 14108 9897 14136 10134
rect 14186 10095 14242 10104
rect 14292 10010 14320 10367
rect 14200 9982 14320 10010
rect 14094 9888 14150 9897
rect 14094 9823 14150 9832
rect 14200 9674 14228 9982
rect 14384 9926 14412 10526
rect 14280 9920 14332 9926
rect 14278 9888 14280 9897
rect 14372 9920 14424 9926
rect 14332 9888 14334 9897
rect 14372 9862 14424 9868
rect 14278 9823 14334 9832
rect 14200 9646 14412 9674
rect 14186 9208 14242 9217
rect 14186 9143 14242 9152
rect 14002 9072 14058 9081
rect 14002 9007 14058 9016
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13910 8120 13966 8129
rect 13910 8055 13966 8064
rect 13912 7948 13964 7954
rect 13832 7908 13912 7936
rect 13912 7890 13964 7896
rect 13818 7848 13874 7857
rect 13728 7812 13780 7818
rect 13818 7783 13874 7792
rect 13728 7754 13780 7760
rect 13740 5778 13768 7754
rect 13832 6662 13860 7783
rect 13924 7750 13952 7890
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13910 7576 13966 7585
rect 13910 7511 13912 7520
rect 13964 7511 13966 7520
rect 13912 7482 13964 7488
rect 13910 7304 13966 7313
rect 13910 7239 13966 7248
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13740 5534 13768 5714
rect 13740 5506 13860 5534
rect 13372 4236 13676 4264
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13174 3904 13230 3913
rect 13174 3839 13230 3848
rect 12806 3768 12862 3777
rect 12806 3703 12862 3712
rect 12716 3528 12768 3534
rect 12820 3505 12848 3703
rect 12716 3470 12768 3476
rect 12806 3496 12862 3505
rect 12622 3224 12678 3233
rect 12532 3188 12584 3194
rect 12622 3159 12678 3168
rect 12728 3176 12756 3470
rect 12806 3431 12862 3440
rect 13176 3460 13228 3466
rect 13176 3402 13228 3408
rect 12794 3292 13102 3301
rect 12794 3290 12800 3292
rect 12856 3290 12880 3292
rect 12936 3290 12960 3292
rect 13016 3290 13040 3292
rect 13096 3290 13102 3292
rect 12856 3238 12858 3290
rect 13038 3238 13040 3290
rect 12794 3236 12800 3238
rect 12856 3236 12880 3238
rect 12936 3236 12960 3238
rect 13016 3236 13040 3238
rect 13096 3236 13102 3238
rect 12794 3227 13102 3236
rect 12728 3148 12940 3176
rect 12532 3130 12584 3136
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12532 3052 12584 3058
rect 12716 3052 12768 3058
rect 12584 3012 12664 3040
rect 12532 2994 12584 3000
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12346 2680 12402 2689
rect 12346 2615 12402 2624
rect 11992 2230 12296 2258
rect 11888 2100 11940 2106
rect 11888 2042 11940 2048
rect 11888 1964 11940 1970
rect 11888 1906 11940 1912
rect 11796 1896 11848 1902
rect 11794 1864 11796 1873
rect 11848 1864 11850 1873
rect 11794 1799 11850 1808
rect 11716 1720 11836 1748
rect 11702 1592 11758 1601
rect 11808 1562 11836 1720
rect 11702 1527 11704 1536
rect 11756 1527 11758 1536
rect 11796 1556 11848 1562
rect 11704 1498 11756 1504
rect 11796 1498 11848 1504
rect 11612 1352 11664 1358
rect 11612 1294 11664 1300
rect 11428 1284 11480 1290
rect 11428 1226 11480 1232
rect 11704 1216 11756 1222
rect 11704 1158 11756 1164
rect 11716 542 11744 1158
rect 11900 649 11928 1906
rect 11886 640 11942 649
rect 11886 575 11942 584
rect 11704 536 11756 542
rect 11704 478 11756 484
rect 11336 468 11388 474
rect 11336 410 11388 416
rect 9864 264 9916 270
rect 9864 206 9916 212
rect 11992 202 12020 2230
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 12084 1834 12112 2042
rect 12164 2032 12216 2038
rect 12164 1974 12216 1980
rect 12176 1834 12204 1974
rect 12360 1970 12388 2615
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12452 2310 12480 2450
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12438 2136 12494 2145
rect 12438 2071 12494 2080
rect 12452 1970 12480 2071
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 12440 1964 12492 1970
rect 12440 1906 12492 1912
rect 12072 1828 12124 1834
rect 12072 1770 12124 1776
rect 12164 1828 12216 1834
rect 12164 1770 12216 1776
rect 12072 1556 12124 1562
rect 12072 1498 12124 1504
rect 12084 1290 12112 1498
rect 12072 1284 12124 1290
rect 12072 1226 12124 1232
rect 12544 1057 12572 2518
rect 12636 2514 12664 3012
rect 12716 2994 12768 3000
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12636 1970 12664 2450
rect 12728 2446 12756 2994
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12728 2020 12756 2382
rect 12820 2310 12848 2858
rect 12912 2310 12940 3148
rect 13188 3074 13216 3402
rect 13096 3058 13216 3074
rect 13084 3052 13216 3058
rect 13136 3046 13216 3052
rect 13268 3052 13320 3058
rect 13084 2994 13136 3000
rect 13268 2994 13320 3000
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 13096 2446 13124 2790
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12900 2304 12952 2310
rect 13004 2292 13032 2382
rect 13004 2281 13216 2292
rect 13004 2272 13230 2281
rect 13004 2264 13174 2272
rect 12900 2246 12952 2252
rect 12794 2204 13102 2213
rect 13174 2207 13230 2216
rect 12794 2202 12800 2204
rect 12856 2202 12880 2204
rect 12936 2202 12960 2204
rect 13016 2202 13040 2204
rect 13096 2202 13102 2204
rect 12856 2150 12858 2202
rect 13038 2150 13040 2202
rect 12794 2148 12800 2150
rect 12856 2148 12880 2150
rect 12936 2148 12960 2150
rect 13016 2148 13040 2150
rect 13096 2148 13102 2150
rect 12794 2139 13102 2148
rect 13280 2122 13308 2994
rect 13188 2094 13308 2122
rect 12808 2032 12860 2038
rect 12728 1992 12808 2020
rect 12808 1974 12860 1980
rect 12624 1964 12676 1970
rect 12624 1906 12676 1912
rect 13084 1896 13136 1902
rect 12990 1864 13046 1873
rect 13188 1884 13216 2094
rect 13268 2032 13320 2038
rect 13268 1974 13320 1980
rect 13136 1856 13216 1884
rect 13084 1838 13136 1844
rect 13280 1816 13308 1974
rect 12990 1799 13046 1808
rect 13004 1766 13032 1799
rect 13188 1788 13308 1816
rect 12992 1760 13044 1766
rect 12992 1702 13044 1708
rect 13188 1494 13216 1788
rect 13266 1728 13322 1737
rect 13266 1663 13322 1672
rect 13280 1562 13308 1663
rect 13268 1556 13320 1562
rect 13268 1498 13320 1504
rect 13176 1488 13228 1494
rect 13176 1430 13228 1436
rect 13268 1352 13320 1358
rect 13188 1300 13268 1306
rect 13188 1294 13320 1300
rect 13084 1284 13136 1290
rect 13188 1278 13308 1294
rect 13188 1272 13216 1278
rect 13136 1244 13216 1272
rect 13084 1226 13136 1232
rect 13268 1216 13320 1222
rect 13268 1158 13320 1164
rect 12794 1116 13102 1125
rect 12794 1114 12800 1116
rect 12856 1114 12880 1116
rect 12936 1114 12960 1116
rect 13016 1114 13040 1116
rect 13096 1114 13102 1116
rect 12856 1062 12858 1114
rect 13038 1062 13040 1114
rect 12794 1060 12800 1062
rect 12856 1060 12880 1062
rect 12936 1060 12960 1062
rect 13016 1060 13040 1062
rect 13096 1060 13102 1062
rect 12530 1048 12586 1057
rect 12794 1051 13102 1060
rect 12530 983 12586 992
rect 13280 513 13308 1158
rect 13372 542 13400 4236
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13464 1834 13492 4014
rect 13556 3126 13584 4082
rect 13740 4049 13768 4150
rect 13726 4040 13782 4049
rect 13726 3975 13782 3984
rect 13726 3904 13782 3913
rect 13726 3839 13782 3848
rect 13740 3466 13768 3839
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13726 3360 13782 3369
rect 13544 3120 13596 3126
rect 13544 3062 13596 3068
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13556 2825 13584 2926
rect 13542 2816 13598 2825
rect 13542 2751 13598 2760
rect 13648 2446 13676 3334
rect 13726 3295 13782 3304
rect 13740 3194 13768 3295
rect 13832 3194 13860 5506
rect 13924 3534 13952 7239
rect 14016 5166 14044 8910
rect 14108 8430 14136 8978
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14094 8120 14150 8129
rect 14094 8055 14150 8064
rect 14108 6186 14136 8055
rect 14200 6798 14228 9143
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14186 6080 14242 6089
rect 14186 6015 14242 6024
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 14108 5012 14136 5646
rect 14016 4984 14136 5012
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13912 3120 13964 3126
rect 13726 3088 13782 3097
rect 13912 3062 13964 3068
rect 13726 3023 13728 3032
rect 13780 3023 13782 3032
rect 13728 2994 13780 3000
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13452 1828 13504 1834
rect 13452 1770 13504 1776
rect 13544 1760 13596 1766
rect 13544 1702 13596 1708
rect 13556 1329 13584 1702
rect 13648 1426 13676 2382
rect 13740 2106 13768 2790
rect 13728 2100 13780 2106
rect 13728 2042 13780 2048
rect 13728 1828 13780 1834
rect 13728 1770 13780 1776
rect 13636 1420 13688 1426
rect 13636 1362 13688 1368
rect 13740 1358 13768 1770
rect 13728 1352 13780 1358
rect 13542 1320 13598 1329
rect 13728 1294 13780 1300
rect 13542 1255 13598 1264
rect 13360 536 13412 542
rect 13266 504 13322 513
rect 13360 478 13412 484
rect 13266 439 13322 448
rect 13832 338 13860 2790
rect 13924 1290 13952 3062
rect 14016 2689 14044 4984
rect 14094 4312 14150 4321
rect 14094 4247 14150 4256
rect 14108 4146 14136 4247
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14108 3913 14136 4082
rect 14094 3904 14150 3913
rect 14094 3839 14150 3848
rect 14096 3120 14148 3126
rect 14094 3088 14096 3097
rect 14148 3088 14150 3097
rect 14094 3023 14150 3032
rect 14002 2680 14058 2689
rect 14200 2650 14228 6015
rect 14292 5030 14320 8978
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14278 4856 14334 4865
rect 14278 4791 14280 4800
rect 14332 4791 14334 4800
rect 14280 4762 14332 4768
rect 14384 4078 14412 9646
rect 14476 5914 14504 12582
rect 14568 11082 14596 13262
rect 14660 12850 14688 14282
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15028 13716 15056 14214
rect 15120 13841 15148 17070
rect 15212 14006 15240 18663
rect 15304 16114 15332 20470
rect 16028 20324 16080 20330
rect 16028 20266 16080 20272
rect 15476 19440 15528 19446
rect 15476 19382 15528 19388
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15106 13832 15162 13841
rect 15304 13784 15332 15914
rect 15106 13767 15162 13776
rect 15212 13756 15332 13784
rect 15028 13688 15148 13716
rect 14768 13628 15076 13637
rect 14768 13626 14774 13628
rect 14830 13626 14854 13628
rect 14910 13626 14934 13628
rect 14990 13626 15014 13628
rect 15070 13626 15076 13628
rect 14830 13574 14832 13626
rect 15012 13574 15014 13626
rect 14768 13572 14774 13574
rect 14830 13572 14854 13574
rect 14910 13572 14934 13574
rect 14990 13572 15014 13574
rect 15070 13572 15076 13574
rect 14768 13563 15076 13572
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14752 12646 14780 13466
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14844 12753 14872 12786
rect 14830 12744 14886 12753
rect 14830 12679 14886 12688
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14768 12540 15076 12549
rect 14768 12538 14774 12540
rect 14830 12538 14854 12540
rect 14910 12538 14934 12540
rect 14990 12538 15014 12540
rect 15070 12538 15076 12540
rect 14830 12486 14832 12538
rect 15012 12486 15014 12538
rect 14768 12484 14774 12486
rect 14830 12484 14854 12486
rect 14910 12484 14934 12486
rect 14990 12484 15014 12486
rect 15070 12484 15076 12486
rect 14768 12475 15076 12484
rect 15120 12442 15148 13688
rect 15212 13530 15240 13756
rect 15290 13696 15346 13705
rect 15290 13631 15346 13640
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15212 12986 15240 13262
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14660 12238 14688 12310
rect 14648 12232 14700 12238
rect 15108 12232 15160 12238
rect 14648 12174 14700 12180
rect 14738 12200 14794 12209
rect 14660 11694 14688 12174
rect 15108 12174 15160 12180
rect 14738 12135 14794 12144
rect 14924 12164 14976 12170
rect 14752 11830 14780 12135
rect 14924 12106 14976 12112
rect 14936 12073 14964 12106
rect 14922 12064 14978 12073
rect 14922 11999 14978 12008
rect 14830 11928 14886 11937
rect 14830 11863 14886 11872
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14844 11540 14872 11863
rect 14660 11512 14872 11540
rect 14660 11150 14688 11512
rect 14768 11452 15076 11461
rect 14768 11450 14774 11452
rect 14830 11450 14854 11452
rect 14910 11450 14934 11452
rect 14990 11450 15014 11452
rect 15070 11450 15076 11452
rect 14830 11398 14832 11450
rect 15012 11398 15014 11450
rect 14768 11396 14774 11398
rect 14830 11396 14854 11398
rect 14910 11396 14934 11398
rect 14990 11396 15014 11398
rect 15070 11396 15076 11398
rect 14768 11387 15076 11396
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 14648 11144 14700 11150
rect 14936 11121 14964 11222
rect 14648 11086 14700 11092
rect 14922 11112 14978 11121
rect 14556 11076 14608 11082
rect 14922 11047 14978 11056
rect 14556 11018 14608 11024
rect 14646 10976 14702 10985
rect 14646 10911 14702 10920
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14568 10198 14596 10678
rect 14660 10606 14688 10911
rect 14830 10840 14886 10849
rect 14830 10775 14886 10784
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14648 10600 14700 10606
rect 14752 10577 14780 10678
rect 14844 10674 14872 10775
rect 15014 10704 15070 10713
rect 14832 10668 14884 10674
rect 15120 10674 15148 12174
rect 15212 11354 15240 12582
rect 15304 11898 15332 13631
rect 15396 13569 15424 17818
rect 15382 13560 15438 13569
rect 15382 13495 15384 13504
rect 15436 13495 15438 13504
rect 15384 13466 15436 13472
rect 15382 13424 15438 13433
rect 15382 13359 15438 13368
rect 15396 12850 15424 13359
rect 15488 12986 15516 19382
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15672 15162 15700 17546
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15474 12880 15530 12889
rect 15384 12844 15436 12850
rect 15474 12815 15530 12824
rect 15384 12786 15436 12792
rect 15396 12617 15424 12786
rect 15382 12608 15438 12617
rect 15382 12543 15438 12552
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15304 11257 15332 11698
rect 15290 11248 15346 11257
rect 15290 11183 15346 11192
rect 15304 11150 15332 11183
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15198 10976 15254 10985
rect 15198 10911 15254 10920
rect 15014 10639 15070 10648
rect 15108 10668 15160 10674
rect 14832 10610 14884 10616
rect 14648 10542 14700 10548
rect 14738 10568 14794 10577
rect 14738 10503 14794 10512
rect 14844 10452 14872 10610
rect 15028 10606 15056 10639
rect 15108 10610 15160 10616
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 14660 10424 14872 10452
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 14556 10056 14608 10062
rect 14660 10044 14688 10424
rect 15212 10418 15240 10911
rect 15290 10840 15346 10849
rect 15290 10775 15292 10784
rect 15344 10775 15346 10784
rect 15292 10746 15344 10752
rect 15120 10390 15240 10418
rect 14768 10364 15076 10373
rect 14768 10362 14774 10364
rect 14830 10362 14854 10364
rect 14910 10362 14934 10364
rect 14990 10362 15014 10364
rect 15070 10362 15076 10364
rect 14830 10310 14832 10362
rect 15012 10310 15014 10362
rect 14768 10308 14774 10310
rect 14830 10308 14854 10310
rect 14910 10308 14934 10310
rect 14990 10308 15014 10310
rect 15070 10308 15076 10310
rect 14768 10299 15076 10308
rect 14740 10260 14792 10266
rect 15120 10248 15148 10390
rect 15290 10296 15346 10305
rect 14740 10202 14792 10208
rect 15028 10220 15148 10248
rect 15212 10254 15290 10282
rect 14608 10016 14688 10044
rect 14556 9998 14608 10004
rect 14556 9920 14608 9926
rect 14554 9888 14556 9897
rect 14608 9888 14610 9897
rect 14752 9874 14780 10202
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14554 9823 14610 9832
rect 14660 9846 14780 9874
rect 14830 9888 14886 9897
rect 14660 9432 14688 9846
rect 14830 9823 14886 9832
rect 14844 9722 14872 9823
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14568 9404 14688 9432
rect 14568 9353 14596 9404
rect 14936 9364 14964 9998
rect 14554 9344 14610 9353
rect 14554 9279 14610 9288
rect 14660 9336 14964 9364
rect 15028 9364 15056 10220
rect 15106 10024 15162 10033
rect 15106 9959 15162 9968
rect 15120 9432 15148 9959
rect 15212 9586 15240 10254
rect 15290 10231 15346 10240
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15120 9404 15240 9432
rect 15028 9336 15148 9364
rect 14554 9072 14610 9081
rect 14554 9007 14610 9016
rect 14568 6322 14596 9007
rect 14660 8974 14688 9336
rect 14768 9276 15076 9285
rect 14768 9274 14774 9276
rect 14830 9274 14854 9276
rect 14910 9274 14934 9276
rect 14990 9274 15014 9276
rect 15070 9274 15076 9276
rect 14830 9222 14832 9274
rect 15012 9222 15014 9274
rect 14768 9220 14774 9222
rect 14830 9220 14854 9222
rect 14910 9220 14934 9222
rect 14990 9220 15014 9222
rect 15070 9220 15076 9222
rect 14768 9211 15076 9220
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14738 8800 14794 8809
rect 14738 8735 14794 8744
rect 14752 8634 14780 8735
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14738 8528 14794 8537
rect 14660 7857 14688 8502
rect 14738 8463 14794 8472
rect 14752 8430 14780 8463
rect 14740 8424 14792 8430
rect 14844 8401 14872 8978
rect 15016 8968 15068 8974
rect 15120 8945 15148 9336
rect 15016 8910 15068 8916
rect 15106 8936 15162 8945
rect 14740 8366 14792 8372
rect 14830 8392 14886 8401
rect 14830 8327 14886 8336
rect 15028 8294 15056 8910
rect 15106 8871 15162 8880
rect 15106 8392 15162 8401
rect 15106 8327 15108 8336
rect 15160 8327 15162 8336
rect 15108 8298 15160 8304
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 14768 8188 15076 8197
rect 14768 8186 14774 8188
rect 14830 8186 14854 8188
rect 14910 8186 14934 8188
rect 14990 8186 15014 8188
rect 15070 8186 15076 8188
rect 14830 8134 14832 8186
rect 15012 8134 15014 8186
rect 14768 8132 14774 8134
rect 14830 8132 14854 8134
rect 14910 8132 14934 8134
rect 14990 8132 15014 8134
rect 15070 8132 15076 8134
rect 14768 8123 15076 8132
rect 15120 8072 15148 8298
rect 15028 8044 15148 8072
rect 14740 7880 14792 7886
rect 14646 7848 14702 7857
rect 14740 7822 14792 7828
rect 14646 7783 14702 7792
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 6390 14688 7686
rect 14752 7478 14780 7822
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14844 7410 14872 7686
rect 15028 7478 15056 8044
rect 15106 7984 15162 7993
rect 15106 7919 15162 7928
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14768 7100 15076 7109
rect 14768 7098 14774 7100
rect 14830 7098 14854 7100
rect 14910 7098 14934 7100
rect 14990 7098 15014 7100
rect 15070 7098 15076 7100
rect 14830 7046 14832 7098
rect 15012 7046 15014 7098
rect 14768 7044 14774 7046
rect 14830 7044 14854 7046
rect 14910 7044 14934 7046
rect 14990 7044 15014 7046
rect 15070 7044 15076 7046
rect 14768 7035 15076 7044
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14752 6798 14780 6938
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14462 5808 14518 5817
rect 14462 5743 14518 5752
rect 14556 5772 14608 5778
rect 14476 5137 14504 5743
rect 14556 5714 14608 5720
rect 14462 5128 14518 5137
rect 14462 5063 14518 5072
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14476 4282 14504 4422
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14370 3904 14426 3913
rect 14292 3738 14320 3878
rect 14370 3839 14426 3848
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14002 2615 14058 2624
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14004 2032 14056 2038
rect 14004 1974 14056 1980
rect 13912 1284 13964 1290
rect 13912 1226 13964 1232
rect 14016 950 14044 1974
rect 14096 1896 14148 1902
rect 14096 1838 14148 1844
rect 14108 1290 14136 1838
rect 14200 1562 14228 2382
rect 14188 1556 14240 1562
rect 14188 1498 14240 1504
rect 14096 1284 14148 1290
rect 14096 1226 14148 1232
rect 14004 944 14056 950
rect 14004 886 14056 892
rect 14108 785 14136 1226
rect 14200 921 14228 1498
rect 14292 1358 14320 3674
rect 14384 3058 14412 3839
rect 14476 3466 14504 4082
rect 14568 3942 14596 5714
rect 14660 4554 14688 6326
rect 14768 6012 15076 6021
rect 14768 6010 14774 6012
rect 14830 6010 14854 6012
rect 14910 6010 14934 6012
rect 14990 6010 15014 6012
rect 15070 6010 15076 6012
rect 14830 5958 14832 6010
rect 15012 5958 15014 6010
rect 14768 5956 14774 5958
rect 14830 5956 14854 5958
rect 14910 5956 14934 5958
rect 14990 5956 15014 5958
rect 15070 5956 15076 5958
rect 14768 5947 15076 5956
rect 15120 5914 15148 7919
rect 15212 6934 15240 9404
rect 15304 8362 15332 9658
rect 15396 8945 15424 12378
rect 15488 12238 15516 12815
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15488 10713 15516 12174
rect 15580 12170 15608 14962
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15672 13297 15700 14826
rect 15658 13288 15714 13297
rect 15658 13223 15714 13232
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15672 12434 15700 12922
rect 15764 12646 15792 17206
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15672 12406 15792 12434
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15672 12209 15700 12310
rect 15658 12200 15714 12209
rect 15568 12164 15620 12170
rect 15658 12135 15714 12144
rect 15568 12106 15620 12112
rect 15474 10704 15530 10713
rect 15474 10639 15530 10648
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15488 10266 15516 10474
rect 15672 10441 15700 10474
rect 15658 10432 15714 10441
rect 15658 10367 15714 10376
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15566 10160 15622 10169
rect 15476 10124 15528 10130
rect 15566 10095 15622 10104
rect 15476 10066 15528 10072
rect 15382 8936 15438 8945
rect 15382 8871 15438 8880
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15396 7886 15424 8774
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15396 7410 15424 7482
rect 15384 7404 15436 7410
rect 15304 7364 15384 7392
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15212 5953 15240 6734
rect 15198 5944 15254 5953
rect 15108 5908 15160 5914
rect 15198 5879 15254 5888
rect 15108 5850 15160 5856
rect 15304 5794 15332 7364
rect 15384 7346 15436 7352
rect 15488 6882 15516 10066
rect 15580 9568 15608 10095
rect 15672 9761 15700 10202
rect 15764 9994 15792 12406
rect 15752 9988 15804 9994
rect 15752 9930 15804 9936
rect 15658 9752 15714 9761
rect 15658 9687 15714 9696
rect 15660 9580 15712 9586
rect 15580 9540 15660 9568
rect 15712 9540 15792 9568
rect 15660 9522 15712 9528
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15580 7274 15608 9114
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15396 6854 15516 6882
rect 15566 6896 15622 6905
rect 15396 6361 15424 6854
rect 15566 6831 15622 6840
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15382 6352 15438 6361
rect 15382 6287 15438 6296
rect 15120 5766 15332 5794
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 14768 4924 15076 4933
rect 14768 4922 14774 4924
rect 14830 4922 14854 4924
rect 14910 4922 14934 4924
rect 14990 4922 15014 4924
rect 15070 4922 15076 4924
rect 14830 4870 14832 4922
rect 15012 4870 15014 4922
rect 14768 4868 14774 4870
rect 14830 4868 14854 4870
rect 14910 4868 14934 4870
rect 14990 4868 15014 4870
rect 15070 4868 15076 4870
rect 14768 4859 15076 4868
rect 15120 4808 15148 5766
rect 15290 5128 15346 5137
rect 15290 5063 15346 5072
rect 15304 5030 15332 5063
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15028 4780 15148 4808
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 14648 4548 14700 4554
rect 14648 4490 14700 4496
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 14646 4448 14702 4457
rect 14646 4383 14702 4392
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14556 3732 14608 3738
rect 14660 3720 14688 4383
rect 14752 4010 14780 4490
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14844 4146 14872 4218
rect 14936 4214 14964 4694
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 15028 4049 15056 4780
rect 15108 4072 15160 4078
rect 15014 4040 15070 4049
rect 14740 4004 14792 4010
rect 15108 4014 15160 4020
rect 15014 3975 15070 3984
rect 14740 3946 14792 3952
rect 14768 3836 15076 3845
rect 14768 3834 14774 3836
rect 14830 3834 14854 3836
rect 14910 3834 14934 3836
rect 14990 3834 15014 3836
rect 15070 3834 15076 3836
rect 14830 3782 14832 3834
rect 15012 3782 15014 3834
rect 14768 3780 14774 3782
rect 14830 3780 14854 3782
rect 14910 3780 14934 3782
rect 14990 3780 15014 3782
rect 15070 3780 15076 3782
rect 14768 3771 15076 3780
rect 14660 3692 14780 3720
rect 14556 3674 14608 3680
rect 14568 3618 14596 3674
rect 14568 3590 14688 3618
rect 14554 3496 14610 3505
rect 14464 3460 14516 3466
rect 14554 3431 14610 3440
rect 14464 3402 14516 3408
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14384 1465 14412 2994
rect 14476 2774 14504 3402
rect 14568 3058 14596 3431
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14660 2854 14688 3590
rect 14752 2990 14780 3692
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 15120 2922 15148 4014
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14476 2746 14596 2774
rect 14464 2032 14516 2038
rect 14568 2009 14596 2746
rect 14660 2417 14688 2790
rect 14768 2748 15076 2757
rect 14768 2746 14774 2748
rect 14830 2746 14854 2748
rect 14910 2746 14934 2748
rect 14990 2746 15014 2748
rect 15070 2746 15076 2748
rect 14830 2694 14832 2746
rect 15012 2694 15014 2746
rect 14768 2692 14774 2694
rect 14830 2692 14854 2694
rect 14910 2692 14934 2694
rect 14990 2692 15014 2694
rect 15070 2692 15076 2694
rect 14768 2683 15076 2692
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 14936 2446 14964 2518
rect 15212 2446 15240 4966
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15304 2961 15332 3878
rect 15396 3058 15424 5782
rect 15488 5370 15516 6734
rect 15580 6662 15608 6831
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15488 3194 15516 4966
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15290 2952 15346 2961
rect 15396 2938 15424 2994
rect 15396 2910 15516 2938
rect 15290 2887 15346 2896
rect 14924 2440 14976 2446
rect 14646 2408 14702 2417
rect 15200 2440 15252 2446
rect 14924 2382 14976 2388
rect 15014 2408 15070 2417
rect 14646 2343 14702 2352
rect 15200 2382 15252 2388
rect 15014 2343 15070 2352
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14844 2145 14872 2246
rect 14830 2136 14886 2145
rect 14830 2071 14886 2080
rect 14464 1974 14516 1980
rect 14554 2000 14610 2009
rect 14476 1562 14504 1974
rect 15028 1970 15056 2343
rect 15488 2106 15516 2910
rect 15580 2650 15608 6054
rect 15672 3233 15700 9318
rect 15764 8974 15792 9540
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15752 8424 15804 8430
rect 15750 8392 15752 8401
rect 15804 8392 15806 8401
rect 15750 8327 15806 8336
rect 15752 7268 15804 7274
rect 15752 7210 15804 7216
rect 15764 5273 15792 7210
rect 15856 5710 15884 15438
rect 15936 15088 15988 15094
rect 15936 15030 15988 15036
rect 15948 12238 15976 15030
rect 16040 13326 16068 20266
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15948 9722 15976 12038
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15750 5264 15806 5273
rect 15856 5234 15884 5646
rect 15750 5199 15806 5208
rect 15844 5228 15896 5234
rect 15764 3670 15792 5199
rect 15844 5170 15896 5176
rect 15752 3664 15804 3670
rect 15752 3606 15804 3612
rect 15658 3224 15714 3233
rect 15658 3159 15714 3168
rect 15750 3088 15806 3097
rect 15856 3058 15884 5170
rect 15948 4826 15976 9046
rect 16040 5642 16068 13262
rect 16132 11558 16160 13670
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16132 10810 16160 11290
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16028 5636 16080 5642
rect 16028 5578 16080 5584
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15948 4214 15976 4762
rect 15936 4208 15988 4214
rect 15936 4150 15988 4156
rect 16026 4176 16082 4185
rect 16026 4111 16028 4120
rect 16080 4111 16082 4120
rect 16028 4082 16080 4088
rect 15750 3023 15806 3032
rect 15844 3052 15896 3058
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 15764 2446 15792 3023
rect 15844 2994 15896 3000
rect 16040 2553 16068 4082
rect 16132 3534 16160 10746
rect 16224 10130 16252 18226
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16316 12782 16344 13738
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16408 12434 16436 13126
rect 16316 12406 16436 12434
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16224 7886 16252 8910
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16224 7290 16252 7822
rect 16316 7449 16344 12406
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 10266 16436 12038
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16408 9489 16436 9930
rect 16394 9480 16450 9489
rect 16394 9415 16450 9424
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16408 7750 16436 8434
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16302 7440 16358 7449
rect 16302 7375 16358 7384
rect 16224 7262 16344 7290
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16224 2650 16252 7142
rect 16316 7002 16344 7262
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16302 6896 16358 6905
rect 16302 6831 16358 6840
rect 16316 3398 16344 6831
rect 16500 3738 16528 16050
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16500 2582 16528 3130
rect 16488 2576 16540 2582
rect 16026 2544 16082 2553
rect 16488 2518 16540 2524
rect 16592 2514 16620 16730
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16684 7818 16712 15302
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16672 6928 16724 6934
rect 16672 6870 16724 6876
rect 16026 2479 16082 2488
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15476 2100 15528 2106
rect 15476 2042 15528 2048
rect 14554 1935 14610 1944
rect 15016 1964 15068 1970
rect 15016 1906 15068 1912
rect 14768 1660 15076 1669
rect 14768 1658 14774 1660
rect 14830 1658 14854 1660
rect 14910 1658 14934 1660
rect 14990 1658 15014 1660
rect 15070 1658 15076 1660
rect 14830 1606 14832 1658
rect 15012 1606 15014 1658
rect 14768 1604 14774 1606
rect 14830 1604 14854 1606
rect 14910 1604 14934 1606
rect 14990 1604 15014 1606
rect 15070 1604 15076 1606
rect 14768 1595 15076 1604
rect 14464 1556 14516 1562
rect 14464 1498 14516 1504
rect 14370 1456 14426 1465
rect 14370 1391 14426 1400
rect 14280 1352 14332 1358
rect 14280 1294 14332 1300
rect 14476 1018 14504 1498
rect 15844 1352 15896 1358
rect 15844 1294 15896 1300
rect 15660 1216 15712 1222
rect 15660 1158 15712 1164
rect 14464 1012 14516 1018
rect 14464 954 14516 960
rect 14186 912 14242 921
rect 14186 847 14242 856
rect 14094 776 14150 785
rect 14094 711 14150 720
rect 13820 332 13872 338
rect 13820 274 13872 280
rect 11980 196 12032 202
rect 11980 138 12032 144
rect 15672 66 15700 1158
rect 15856 814 15884 1294
rect 15844 808 15896 814
rect 15844 750 15896 756
rect 16040 406 16068 2382
rect 16684 882 16712 6870
rect 16776 4282 16804 17002
rect 16868 11354 16896 18634
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16868 10470 16896 11154
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16764 4276 16816 4282
rect 16764 4218 16816 4224
rect 16868 4078 16896 9998
rect 16960 7546 16988 22374
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 17052 2774 17080 18702
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17144 6322 17172 18022
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17236 4321 17264 19994
rect 17222 4312 17278 4321
rect 17222 4247 17278 4256
rect 16868 2746 17080 2774
rect 16672 876 16724 882
rect 16672 818 16724 824
rect 16868 678 16896 2746
rect 17328 1766 17356 20402
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17316 1760 17368 1766
rect 17316 1702 17368 1708
rect 17420 1562 17448 20198
rect 17592 19236 17644 19242
rect 17592 19178 17644 19184
rect 17498 13152 17554 13161
rect 17498 13087 17554 13096
rect 17512 6390 17540 13087
rect 17500 6384 17552 6390
rect 17500 6326 17552 6332
rect 17604 3369 17632 19178
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17696 6769 17724 8230
rect 17682 6760 17738 6769
rect 17682 6695 17738 6704
rect 17590 3360 17646 3369
rect 17590 3295 17646 3304
rect 17408 1556 17460 1562
rect 17408 1498 17460 1504
rect 16856 672 16908 678
rect 16856 614 16908 620
rect 16028 400 16080 406
rect 16028 342 16080 348
rect 7748 60 7800 66
rect 7748 2 7800 8
rect 15660 60 15712 66
rect 15660 2 15712 8
<< via2 >>
rect 1582 23160 1638 23216
rect 1490 22500 1546 22536
rect 1490 22480 1492 22500
rect 1492 22480 1544 22500
rect 1544 22480 1546 22500
rect 4904 22874 4960 22876
rect 4984 22874 5040 22876
rect 5064 22874 5120 22876
rect 5144 22874 5200 22876
rect 4904 22822 4950 22874
rect 4950 22822 4960 22874
rect 4984 22822 5014 22874
rect 5014 22822 5026 22874
rect 5026 22822 5040 22874
rect 5064 22822 5078 22874
rect 5078 22822 5090 22874
rect 5090 22822 5120 22874
rect 5144 22822 5154 22874
rect 5154 22822 5200 22874
rect 4904 22820 4960 22822
rect 4984 22820 5040 22822
rect 5064 22820 5120 22822
rect 5144 22820 5200 22822
rect 8852 22874 8908 22876
rect 8932 22874 8988 22876
rect 9012 22874 9068 22876
rect 9092 22874 9148 22876
rect 8852 22822 8898 22874
rect 8898 22822 8908 22874
rect 8932 22822 8962 22874
rect 8962 22822 8974 22874
rect 8974 22822 8988 22874
rect 9012 22822 9026 22874
rect 9026 22822 9038 22874
rect 9038 22822 9068 22874
rect 9092 22822 9102 22874
rect 9102 22822 9148 22874
rect 8852 22820 8908 22822
rect 8932 22820 8988 22822
rect 9012 22820 9068 22822
rect 9092 22820 9148 22822
rect 12800 22874 12856 22876
rect 12880 22874 12936 22876
rect 12960 22874 13016 22876
rect 13040 22874 13096 22876
rect 12800 22822 12846 22874
rect 12846 22822 12856 22874
rect 12880 22822 12910 22874
rect 12910 22822 12922 22874
rect 12922 22822 12936 22874
rect 12960 22822 12974 22874
rect 12974 22822 12986 22874
rect 12986 22822 13016 22874
rect 13040 22822 13050 22874
rect 13050 22822 13096 22874
rect 12800 22820 12856 22822
rect 12880 22820 12936 22822
rect 12960 22820 13016 22822
rect 13040 22820 13096 22822
rect 2930 22330 2986 22332
rect 3010 22330 3066 22332
rect 3090 22330 3146 22332
rect 3170 22330 3226 22332
rect 2930 22278 2976 22330
rect 2976 22278 2986 22330
rect 3010 22278 3040 22330
rect 3040 22278 3052 22330
rect 3052 22278 3066 22330
rect 3090 22278 3104 22330
rect 3104 22278 3116 22330
rect 3116 22278 3146 22330
rect 3170 22278 3180 22330
rect 3180 22278 3226 22330
rect 2930 22276 2986 22278
rect 3010 22276 3066 22278
rect 3090 22276 3146 22278
rect 3170 22276 3226 22278
rect 6878 22330 6934 22332
rect 6958 22330 7014 22332
rect 7038 22330 7094 22332
rect 7118 22330 7174 22332
rect 6878 22278 6924 22330
rect 6924 22278 6934 22330
rect 6958 22278 6988 22330
rect 6988 22278 7000 22330
rect 7000 22278 7014 22330
rect 7038 22278 7052 22330
rect 7052 22278 7064 22330
rect 7064 22278 7094 22330
rect 7118 22278 7128 22330
rect 7128 22278 7174 22330
rect 6878 22276 6934 22278
rect 6958 22276 7014 22278
rect 7038 22276 7094 22278
rect 7118 22276 7174 22278
rect 10826 22330 10882 22332
rect 10906 22330 10962 22332
rect 10986 22330 11042 22332
rect 11066 22330 11122 22332
rect 10826 22278 10872 22330
rect 10872 22278 10882 22330
rect 10906 22278 10936 22330
rect 10936 22278 10948 22330
rect 10948 22278 10962 22330
rect 10986 22278 11000 22330
rect 11000 22278 11012 22330
rect 11012 22278 11042 22330
rect 11066 22278 11076 22330
rect 11076 22278 11122 22330
rect 10826 22276 10882 22278
rect 10906 22276 10962 22278
rect 10986 22276 11042 22278
rect 11066 22276 11122 22278
rect 2410 21664 2466 21720
rect 18 17720 74 17776
rect 478 19216 534 19272
rect 938 17584 994 17640
rect 570 16224 626 16280
rect 478 8200 534 8256
rect 18 2488 74 2544
rect 662 15408 718 15464
rect 754 13776 810 13832
rect 1030 2896 1086 2952
rect 14774 22330 14830 22332
rect 14854 22330 14910 22332
rect 14934 22330 14990 22332
rect 15014 22330 15070 22332
rect 14774 22278 14820 22330
rect 14820 22278 14830 22330
rect 14854 22278 14884 22330
rect 14884 22278 14896 22330
rect 14896 22278 14910 22330
rect 14934 22278 14948 22330
rect 14948 22278 14960 22330
rect 14960 22278 14990 22330
rect 15014 22278 15024 22330
rect 15024 22278 15070 22330
rect 14774 22276 14830 22278
rect 14854 22276 14910 22278
rect 14934 22276 14990 22278
rect 15014 22276 15070 22278
rect 2930 21242 2986 21244
rect 3010 21242 3066 21244
rect 3090 21242 3146 21244
rect 3170 21242 3226 21244
rect 2930 21190 2976 21242
rect 2976 21190 2986 21242
rect 3010 21190 3040 21242
rect 3040 21190 3052 21242
rect 3052 21190 3066 21242
rect 3090 21190 3104 21242
rect 3104 21190 3116 21242
rect 3116 21190 3146 21242
rect 3170 21190 3180 21242
rect 3180 21190 3226 21242
rect 2930 21188 2986 21190
rect 3010 21188 3066 21190
rect 3090 21188 3146 21190
rect 3170 21188 3226 21190
rect 1398 15680 1454 15736
rect 1490 14184 1546 14240
rect 1582 13368 1638 13424
rect 1582 12960 1638 13016
rect 1950 16360 2006 16416
rect 1858 13388 1914 13424
rect 1858 13368 1860 13388
rect 1860 13368 1912 13388
rect 1912 13368 1914 13388
rect 2226 15952 2282 16008
rect 3146 20304 3202 20360
rect 2778 20168 2834 20224
rect 2930 20154 2986 20156
rect 3010 20154 3066 20156
rect 3090 20154 3146 20156
rect 3170 20154 3226 20156
rect 2930 20102 2976 20154
rect 2976 20102 2986 20154
rect 3010 20102 3040 20154
rect 3040 20102 3052 20154
rect 3052 20102 3066 20154
rect 3090 20102 3104 20154
rect 3104 20102 3116 20154
rect 3116 20102 3146 20154
rect 3170 20102 3180 20154
rect 3180 20102 3226 20154
rect 2930 20100 2986 20102
rect 3010 20100 3066 20102
rect 3090 20100 3146 20102
rect 3170 20100 3226 20102
rect 3146 19896 3202 19952
rect 2870 19780 2926 19816
rect 2870 19760 2872 19780
rect 2872 19760 2924 19780
rect 2924 19760 2926 19780
rect 2594 19388 2596 19408
rect 2596 19388 2648 19408
rect 2648 19388 2650 19408
rect 2594 19352 2650 19388
rect 2594 18808 2650 18864
rect 3330 19624 3386 19680
rect 3330 19216 3386 19272
rect 2930 19066 2986 19068
rect 3010 19066 3066 19068
rect 3090 19066 3146 19068
rect 3170 19066 3226 19068
rect 2930 19014 2976 19066
rect 2976 19014 2986 19066
rect 3010 19014 3040 19066
rect 3040 19014 3052 19066
rect 3052 19014 3066 19066
rect 3090 19014 3104 19066
rect 3104 19014 3116 19066
rect 3116 19014 3146 19066
rect 3170 19014 3180 19066
rect 3180 19014 3226 19066
rect 2930 19012 2986 19014
rect 3010 19012 3066 19014
rect 3090 19012 3146 19014
rect 3170 19012 3226 19014
rect 2410 16496 2466 16552
rect 2410 16360 2466 16416
rect 2686 18128 2742 18184
rect 2686 16496 2742 16552
rect 2410 13232 2466 13288
rect 2226 12824 2282 12880
rect 1950 12688 2006 12744
rect 1766 10668 1822 10704
rect 1766 10648 1768 10668
rect 1768 10648 1820 10668
rect 1820 10648 1822 10668
rect 1490 3168 1546 3224
rect 1306 1400 1362 1456
rect 2594 14592 2650 14648
rect 2410 12144 2466 12200
rect 2318 12008 2374 12064
rect 2226 11736 2282 11792
rect 2226 10512 2282 10568
rect 2134 9460 2136 9480
rect 2136 9460 2188 9480
rect 2188 9460 2190 9480
rect 2134 9424 2190 9460
rect 1490 1264 1546 1320
rect 2318 6160 2374 6216
rect 2594 12280 2650 12336
rect 2594 11872 2650 11928
rect 3054 18536 3110 18592
rect 3606 20168 3662 20224
rect 2930 17978 2986 17980
rect 3010 17978 3066 17980
rect 3090 17978 3146 17980
rect 3170 17978 3226 17980
rect 2930 17926 2976 17978
rect 2976 17926 2986 17978
rect 3010 17926 3040 17978
rect 3040 17926 3052 17978
rect 3052 17926 3066 17978
rect 3090 17926 3104 17978
rect 3104 17926 3116 17978
rect 3116 17926 3146 17978
rect 3170 17926 3180 17978
rect 3180 17926 3226 17978
rect 2930 17924 2986 17926
rect 3010 17924 3066 17926
rect 3090 17924 3146 17926
rect 3170 17924 3226 17926
rect 3330 17176 3386 17232
rect 2930 16890 2986 16892
rect 3010 16890 3066 16892
rect 3090 16890 3146 16892
rect 3170 16890 3226 16892
rect 2930 16838 2976 16890
rect 2976 16838 2986 16890
rect 3010 16838 3040 16890
rect 3040 16838 3052 16890
rect 3052 16838 3066 16890
rect 3090 16838 3104 16890
rect 3104 16838 3116 16890
rect 3116 16838 3146 16890
rect 3170 16838 3180 16890
rect 3180 16838 3226 16890
rect 2930 16836 2986 16838
rect 3010 16836 3066 16838
rect 3090 16836 3146 16838
rect 3170 16836 3226 16838
rect 2930 15802 2986 15804
rect 3010 15802 3066 15804
rect 3090 15802 3146 15804
rect 3170 15802 3226 15804
rect 2930 15750 2976 15802
rect 2976 15750 2986 15802
rect 3010 15750 3040 15802
rect 3040 15750 3052 15802
rect 3052 15750 3066 15802
rect 3090 15750 3104 15802
rect 3104 15750 3116 15802
rect 3116 15750 3146 15802
rect 3170 15750 3180 15802
rect 3180 15750 3226 15802
rect 2930 15748 2986 15750
rect 3010 15748 3066 15750
rect 3090 15748 3146 15750
rect 3170 15748 3226 15750
rect 2930 14714 2986 14716
rect 3010 14714 3066 14716
rect 3090 14714 3146 14716
rect 3170 14714 3226 14716
rect 2930 14662 2976 14714
rect 2976 14662 2986 14714
rect 3010 14662 3040 14714
rect 3040 14662 3052 14714
rect 3052 14662 3066 14714
rect 3090 14662 3104 14714
rect 3104 14662 3116 14714
rect 3116 14662 3146 14714
rect 3170 14662 3180 14714
rect 3180 14662 3226 14714
rect 2930 14660 2986 14662
rect 3010 14660 3066 14662
rect 3090 14660 3146 14662
rect 3170 14660 3226 14662
rect 2962 13812 2964 13832
rect 2964 13812 3016 13832
rect 3016 13812 3018 13832
rect 2962 13776 3018 13812
rect 2930 13626 2986 13628
rect 3010 13626 3066 13628
rect 3090 13626 3146 13628
rect 3170 13626 3226 13628
rect 2930 13574 2976 13626
rect 2976 13574 2986 13626
rect 3010 13574 3040 13626
rect 3040 13574 3052 13626
rect 3052 13574 3066 13626
rect 3090 13574 3104 13626
rect 3104 13574 3116 13626
rect 3116 13574 3146 13626
rect 3170 13574 3180 13626
rect 3180 13574 3226 13626
rect 2930 13572 2986 13574
rect 3010 13572 3066 13574
rect 3090 13572 3146 13574
rect 3170 13572 3226 13574
rect 2870 13404 2872 13424
rect 2872 13404 2924 13424
rect 2924 13404 2926 13424
rect 2870 13368 2926 13404
rect 3146 13368 3202 13424
rect 2930 12538 2986 12540
rect 3010 12538 3066 12540
rect 3090 12538 3146 12540
rect 3170 12538 3226 12540
rect 2930 12486 2976 12538
rect 2976 12486 2986 12538
rect 3010 12486 3040 12538
rect 3040 12486 3052 12538
rect 3052 12486 3066 12538
rect 3090 12486 3104 12538
rect 3104 12486 3116 12538
rect 3116 12486 3146 12538
rect 3170 12486 3180 12538
rect 3180 12486 3226 12538
rect 2930 12484 2986 12486
rect 3010 12484 3066 12486
rect 3090 12484 3146 12486
rect 3170 12484 3226 12486
rect 2594 10784 2650 10840
rect 3146 11872 3202 11928
rect 3422 12180 3424 12200
rect 3424 12180 3476 12200
rect 3476 12180 3478 12200
rect 3422 12144 3478 12180
rect 3422 12008 3478 12064
rect 3790 20032 3846 20088
rect 3698 18672 3754 18728
rect 4904 21786 4960 21788
rect 4984 21786 5040 21788
rect 5064 21786 5120 21788
rect 5144 21786 5200 21788
rect 4904 21734 4950 21786
rect 4950 21734 4960 21786
rect 4984 21734 5014 21786
rect 5014 21734 5026 21786
rect 5026 21734 5040 21786
rect 5064 21734 5078 21786
rect 5078 21734 5090 21786
rect 5090 21734 5120 21786
rect 5144 21734 5154 21786
rect 5154 21734 5200 21786
rect 4904 21732 4960 21734
rect 4984 21732 5040 21734
rect 5064 21732 5120 21734
rect 5144 21732 5200 21734
rect 3974 19896 4030 19952
rect 4904 20698 4960 20700
rect 4984 20698 5040 20700
rect 5064 20698 5120 20700
rect 5144 20698 5200 20700
rect 4904 20646 4950 20698
rect 4950 20646 4960 20698
rect 4984 20646 5014 20698
rect 5014 20646 5026 20698
rect 5026 20646 5040 20698
rect 5064 20646 5078 20698
rect 5078 20646 5090 20698
rect 5090 20646 5120 20698
rect 5144 20646 5154 20698
rect 5154 20646 5200 20698
rect 4904 20644 4960 20646
rect 4984 20644 5040 20646
rect 5064 20644 5120 20646
rect 5144 20644 5200 20646
rect 3790 18400 3846 18456
rect 4066 18808 4122 18864
rect 4066 18128 4122 18184
rect 4066 18028 4068 18048
rect 4068 18028 4120 18048
rect 4120 18028 4122 18048
rect 4066 17992 4122 18028
rect 3974 15952 4030 16008
rect 4066 14184 4122 14240
rect 3974 13932 4030 13968
rect 3974 13912 3976 13932
rect 3976 13912 4028 13932
rect 4028 13912 4030 13932
rect 3882 13504 3938 13560
rect 3882 13096 3938 13152
rect 3698 12688 3754 12744
rect 3606 12552 3662 12608
rect 2930 11450 2986 11452
rect 3010 11450 3066 11452
rect 3090 11450 3146 11452
rect 3170 11450 3226 11452
rect 2930 11398 2976 11450
rect 2976 11398 2986 11450
rect 3010 11398 3040 11450
rect 3040 11398 3052 11450
rect 3052 11398 3066 11450
rect 3090 11398 3104 11450
rect 3104 11398 3116 11450
rect 3116 11398 3146 11450
rect 3170 11398 3180 11450
rect 3180 11398 3226 11450
rect 2930 11396 2986 11398
rect 3010 11396 3066 11398
rect 3090 11396 3146 11398
rect 3170 11396 3226 11398
rect 2962 11212 3018 11248
rect 2962 11192 2964 11212
rect 2964 11192 3016 11212
rect 3016 11192 3018 11212
rect 3606 11328 3662 11384
rect 2870 11056 2926 11112
rect 2930 10362 2986 10364
rect 3010 10362 3066 10364
rect 3090 10362 3146 10364
rect 3170 10362 3226 10364
rect 2930 10310 2976 10362
rect 2976 10310 2986 10362
rect 3010 10310 3040 10362
rect 3040 10310 3052 10362
rect 3052 10310 3066 10362
rect 3090 10310 3104 10362
rect 3104 10310 3116 10362
rect 3116 10310 3146 10362
rect 3170 10310 3180 10362
rect 3180 10310 3226 10362
rect 2930 10308 2986 10310
rect 3010 10308 3066 10310
rect 3090 10308 3146 10310
rect 3170 10308 3226 10310
rect 3146 10124 3202 10160
rect 3146 10104 3148 10124
rect 3148 10104 3200 10124
rect 3200 10104 3202 10124
rect 3146 9968 3202 10024
rect 2686 8608 2742 8664
rect 2686 6840 2742 6896
rect 2930 9274 2986 9276
rect 3010 9274 3066 9276
rect 3090 9274 3146 9276
rect 3170 9274 3226 9276
rect 2930 9222 2976 9274
rect 2976 9222 2986 9274
rect 3010 9222 3040 9274
rect 3040 9222 3052 9274
rect 3052 9222 3066 9274
rect 3090 9222 3104 9274
rect 3104 9222 3116 9274
rect 3116 9222 3146 9274
rect 3170 9222 3180 9274
rect 3180 9222 3226 9274
rect 2930 9220 2986 9222
rect 3010 9220 3066 9222
rect 3090 9220 3146 9222
rect 3170 9220 3226 9222
rect 2930 8186 2986 8188
rect 3010 8186 3066 8188
rect 3090 8186 3146 8188
rect 3170 8186 3226 8188
rect 2930 8134 2976 8186
rect 2976 8134 2986 8186
rect 3010 8134 3040 8186
rect 3040 8134 3052 8186
rect 3052 8134 3066 8186
rect 3090 8134 3104 8186
rect 3104 8134 3116 8186
rect 3116 8134 3146 8186
rect 3170 8134 3180 8186
rect 3180 8134 3226 8186
rect 2930 8132 2986 8134
rect 3010 8132 3066 8134
rect 3090 8132 3146 8134
rect 3170 8132 3226 8134
rect 2930 7098 2986 7100
rect 3010 7098 3066 7100
rect 3090 7098 3146 7100
rect 3170 7098 3226 7100
rect 2930 7046 2976 7098
rect 2976 7046 2986 7098
rect 3010 7046 3040 7098
rect 3040 7046 3052 7098
rect 3052 7046 3066 7098
rect 3090 7046 3104 7098
rect 3104 7046 3116 7098
rect 3116 7046 3146 7098
rect 3170 7046 3180 7098
rect 3180 7046 3226 7098
rect 2930 7044 2986 7046
rect 3010 7044 3066 7046
rect 3090 7044 3146 7046
rect 3170 7044 3226 7046
rect 2686 5752 2742 5808
rect 2502 4664 2558 4720
rect 1950 584 2006 640
rect 2930 6010 2986 6012
rect 3010 6010 3066 6012
rect 3090 6010 3146 6012
rect 3170 6010 3226 6012
rect 2930 5958 2976 6010
rect 2976 5958 2986 6010
rect 3010 5958 3040 6010
rect 3040 5958 3052 6010
rect 3052 5958 3066 6010
rect 3090 5958 3104 6010
rect 3104 5958 3116 6010
rect 3116 5958 3146 6010
rect 3170 5958 3180 6010
rect 3180 5958 3226 6010
rect 2930 5956 2986 5958
rect 3010 5956 3066 5958
rect 3090 5956 3146 5958
rect 3170 5956 3226 5958
rect 2778 5208 2834 5264
rect 3330 4936 3386 4992
rect 2930 4922 2986 4924
rect 3010 4922 3066 4924
rect 3090 4922 3146 4924
rect 3170 4922 3226 4924
rect 2930 4870 2976 4922
rect 2976 4870 2986 4922
rect 3010 4870 3040 4922
rect 3040 4870 3052 4922
rect 3052 4870 3066 4922
rect 3090 4870 3104 4922
rect 3104 4870 3116 4922
rect 3116 4870 3146 4922
rect 3170 4870 3180 4922
rect 3180 4870 3226 4922
rect 2930 4868 2986 4870
rect 3010 4868 3066 4870
rect 3090 4868 3146 4870
rect 3170 4868 3226 4870
rect 2870 4256 2926 4312
rect 2930 3834 2986 3836
rect 3010 3834 3066 3836
rect 3090 3834 3146 3836
rect 3170 3834 3226 3836
rect 2930 3782 2976 3834
rect 2976 3782 2986 3834
rect 3010 3782 3040 3834
rect 3040 3782 3052 3834
rect 3052 3782 3066 3834
rect 3090 3782 3104 3834
rect 3104 3782 3116 3834
rect 3116 3782 3146 3834
rect 3170 3782 3180 3834
rect 3180 3782 3226 3834
rect 2930 3780 2986 3782
rect 3010 3780 3066 3782
rect 3090 3780 3146 3782
rect 3170 3780 3226 3782
rect 3146 3476 3148 3496
rect 3148 3476 3200 3496
rect 3200 3476 3202 3496
rect 3146 3440 3202 3476
rect 3514 10376 3570 10432
rect 3606 8492 3662 8528
rect 3606 8472 3608 8492
rect 3608 8472 3660 8492
rect 3660 8472 3662 8492
rect 3606 7248 3662 7304
rect 3514 6840 3570 6896
rect 3882 12164 3938 12200
rect 3882 12144 3884 12164
rect 3884 12144 3936 12164
rect 3936 12144 3938 12164
rect 3882 10920 3938 10976
rect 4066 13096 4122 13152
rect 4342 20304 4398 20360
rect 4342 17176 4398 17232
rect 5814 20204 5816 20224
rect 5816 20204 5868 20224
rect 5868 20204 5870 20224
rect 4710 20032 4766 20088
rect 5538 20032 5594 20088
rect 4710 19624 4766 19680
rect 4904 19610 4960 19612
rect 4984 19610 5040 19612
rect 5064 19610 5120 19612
rect 5144 19610 5200 19612
rect 4904 19558 4950 19610
rect 4950 19558 4960 19610
rect 4984 19558 5014 19610
rect 5014 19558 5026 19610
rect 5026 19558 5040 19610
rect 5064 19558 5078 19610
rect 5078 19558 5090 19610
rect 5090 19558 5120 19610
rect 5144 19558 5154 19610
rect 5154 19558 5200 19610
rect 4904 19556 4960 19558
rect 4984 19556 5040 19558
rect 5064 19556 5120 19558
rect 5144 19556 5200 19558
rect 4710 19352 4766 19408
rect 4710 19216 4766 19272
rect 5262 19388 5264 19408
rect 5264 19388 5316 19408
rect 5316 19388 5318 19408
rect 5262 19352 5318 19388
rect 4710 18400 4766 18456
rect 4526 16360 4582 16416
rect 4618 15272 4674 15328
rect 4526 14592 4582 14648
rect 4434 14320 4490 14376
rect 4904 18522 4960 18524
rect 4984 18522 5040 18524
rect 5064 18522 5120 18524
rect 5144 18522 5200 18524
rect 4904 18470 4950 18522
rect 4950 18470 4960 18522
rect 4984 18470 5014 18522
rect 5014 18470 5026 18522
rect 5026 18470 5040 18522
rect 5064 18470 5078 18522
rect 5078 18470 5090 18522
rect 5090 18470 5120 18522
rect 5144 18470 5154 18522
rect 5154 18470 5200 18522
rect 4904 18468 4960 18470
rect 4984 18468 5040 18470
rect 5064 18468 5120 18470
rect 5144 18468 5200 18470
rect 5170 17584 5226 17640
rect 4904 17434 4960 17436
rect 4984 17434 5040 17436
rect 5064 17434 5120 17436
rect 5144 17434 5200 17436
rect 4904 17382 4950 17434
rect 4950 17382 4960 17434
rect 4984 17382 5014 17434
rect 5014 17382 5026 17434
rect 5026 17382 5040 17434
rect 5064 17382 5078 17434
rect 5078 17382 5090 17434
rect 5090 17382 5120 17434
rect 5144 17382 5154 17434
rect 5154 17382 5200 17434
rect 4904 17380 4960 17382
rect 4984 17380 5040 17382
rect 5064 17380 5120 17382
rect 5144 17380 5200 17382
rect 4802 16496 4858 16552
rect 4904 16346 4960 16348
rect 4984 16346 5040 16348
rect 5064 16346 5120 16348
rect 5144 16346 5200 16348
rect 4904 16294 4950 16346
rect 4950 16294 4960 16346
rect 4984 16294 5014 16346
rect 5014 16294 5026 16346
rect 5026 16294 5040 16346
rect 5064 16294 5078 16346
rect 5078 16294 5090 16346
rect 5090 16294 5120 16346
rect 5144 16294 5154 16346
rect 5154 16294 5200 16346
rect 4904 16292 4960 16294
rect 4984 16292 5040 16294
rect 5064 16292 5120 16294
rect 5144 16292 5200 16294
rect 5078 15816 5134 15872
rect 4904 15258 4960 15260
rect 4984 15258 5040 15260
rect 5064 15258 5120 15260
rect 5144 15258 5200 15260
rect 4904 15206 4950 15258
rect 4950 15206 4960 15258
rect 4984 15206 5014 15258
rect 5014 15206 5026 15258
rect 5026 15206 5040 15258
rect 5064 15206 5078 15258
rect 5078 15206 5090 15258
rect 5090 15206 5120 15258
rect 5144 15206 5154 15258
rect 5154 15206 5200 15258
rect 4904 15204 4960 15206
rect 4984 15204 5040 15206
rect 5064 15204 5120 15206
rect 5144 15204 5200 15206
rect 4894 14864 4950 14920
rect 4802 14456 4858 14512
rect 4526 13388 4582 13424
rect 4526 13368 4528 13388
rect 4528 13368 4580 13388
rect 4580 13368 4582 13388
rect 4526 13232 4582 13288
rect 4342 12552 4398 12608
rect 4066 12008 4122 12064
rect 4066 11756 4122 11792
rect 4066 11736 4068 11756
rect 4068 11736 4120 11756
rect 4120 11736 4122 11756
rect 4250 12144 4306 12200
rect 4526 12416 4582 12472
rect 4434 12144 4490 12200
rect 4158 11464 4214 11520
rect 4066 11328 4122 11384
rect 4250 11212 4306 11248
rect 4250 11192 4252 11212
rect 4252 11192 4304 11212
rect 4304 11192 4306 11212
rect 4434 10648 4490 10704
rect 4066 9716 4122 9752
rect 4066 9696 4068 9716
rect 4068 9696 4120 9716
rect 4120 9696 4122 9716
rect 3698 6296 3754 6352
rect 3606 4256 3662 4312
rect 3790 4564 3792 4584
rect 3792 4564 3844 4584
rect 3844 4564 3846 4584
rect 3790 4528 3846 4564
rect 3698 3576 3754 3632
rect 3882 3576 3938 3632
rect 2930 2746 2986 2748
rect 3010 2746 3066 2748
rect 3090 2746 3146 2748
rect 3170 2746 3226 2748
rect 2930 2694 2976 2746
rect 2976 2694 2986 2746
rect 3010 2694 3040 2746
rect 3040 2694 3052 2746
rect 3052 2694 3066 2746
rect 3090 2694 3104 2746
rect 3104 2694 3116 2746
rect 3116 2694 3146 2746
rect 3170 2694 3180 2746
rect 3180 2694 3226 2746
rect 2930 2692 2986 2694
rect 3010 2692 3066 2694
rect 3090 2692 3146 2694
rect 3170 2692 3226 2694
rect 2870 2488 2926 2544
rect 2502 2352 2558 2408
rect 3146 2352 3202 2408
rect 2686 1844 2688 1864
rect 2688 1844 2740 1864
rect 2740 1844 2742 1864
rect 2686 1808 2742 1844
rect 4342 9560 4398 9616
rect 4066 8472 4122 8528
rect 4434 8608 4490 8664
rect 4066 8372 4068 8392
rect 4068 8372 4120 8392
rect 4120 8372 4122 8392
rect 4066 8336 4122 8372
rect 4066 6160 4122 6216
rect 4066 5652 4068 5672
rect 4068 5652 4120 5672
rect 4120 5652 4122 5672
rect 4066 5616 4122 5652
rect 4342 8472 4398 8528
rect 4158 3304 4214 3360
rect 2930 1658 2986 1660
rect 3010 1658 3066 1660
rect 3090 1658 3146 1660
rect 3170 1658 3226 1660
rect 2930 1606 2976 1658
rect 2976 1606 2986 1658
rect 3010 1606 3040 1658
rect 3040 1606 3052 1658
rect 3052 1606 3066 1658
rect 3090 1606 3104 1658
rect 3104 1606 3116 1658
rect 3116 1606 3146 1658
rect 3170 1606 3180 1658
rect 3180 1606 3226 1658
rect 2930 1604 2986 1606
rect 3010 1604 3066 1606
rect 3090 1604 3146 1606
rect 3170 1604 3226 1606
rect 2962 1300 2964 1320
rect 2964 1300 3016 1320
rect 3016 1300 3018 1320
rect 2962 1264 3018 1300
rect 4158 2352 4214 2408
rect 4066 1536 4122 1592
rect 4434 3848 4490 3904
rect 4710 13676 4712 13696
rect 4712 13676 4764 13696
rect 4764 13676 4766 13696
rect 4710 13640 4766 13676
rect 4710 12980 4766 13016
rect 4710 12960 4712 12980
rect 4712 12960 4764 12980
rect 4764 12960 4766 12980
rect 4904 14170 4960 14172
rect 4984 14170 5040 14172
rect 5064 14170 5120 14172
rect 5144 14170 5200 14172
rect 4904 14118 4950 14170
rect 4950 14118 4960 14170
rect 4984 14118 5014 14170
rect 5014 14118 5026 14170
rect 5026 14118 5040 14170
rect 5064 14118 5078 14170
rect 5078 14118 5090 14170
rect 5090 14118 5120 14170
rect 5144 14118 5154 14170
rect 5154 14118 5200 14170
rect 4904 14116 4960 14118
rect 4984 14116 5040 14118
rect 5064 14116 5120 14118
rect 5144 14116 5200 14118
rect 4894 13776 4950 13832
rect 4894 13232 4950 13288
rect 4904 13082 4960 13084
rect 4984 13082 5040 13084
rect 5064 13082 5120 13084
rect 5144 13082 5200 13084
rect 4904 13030 4950 13082
rect 4950 13030 4960 13082
rect 4984 13030 5014 13082
rect 5014 13030 5026 13082
rect 5026 13030 5040 13082
rect 5064 13030 5078 13082
rect 5078 13030 5090 13082
rect 5090 13030 5120 13082
rect 5144 13030 5154 13082
rect 5154 13030 5200 13082
rect 4904 13028 4960 13030
rect 4984 13028 5040 13030
rect 5064 13028 5120 13030
rect 5144 13028 5200 13030
rect 4894 12688 4950 12744
rect 4802 12416 4858 12472
rect 4986 12300 5042 12336
rect 4986 12280 4988 12300
rect 4988 12280 5040 12300
rect 5040 12280 5042 12300
rect 5170 12552 5226 12608
rect 5078 12144 5134 12200
rect 4904 11994 4960 11996
rect 4984 11994 5040 11996
rect 5064 11994 5120 11996
rect 5144 11994 5200 11996
rect 4904 11942 4950 11994
rect 4950 11942 4960 11994
rect 4984 11942 5014 11994
rect 5014 11942 5026 11994
rect 5026 11942 5040 11994
rect 5064 11942 5078 11994
rect 5078 11942 5090 11994
rect 5090 11942 5120 11994
rect 5144 11942 5154 11994
rect 5154 11942 5200 11994
rect 4904 11940 4960 11942
rect 4984 11940 5040 11942
rect 5064 11940 5120 11942
rect 5144 11940 5200 11942
rect 5170 11756 5226 11792
rect 5170 11736 5172 11756
rect 5172 11736 5224 11756
rect 5224 11736 5226 11756
rect 5078 11464 5134 11520
rect 4802 11328 4858 11384
rect 4710 10920 4766 10976
rect 4710 10512 4766 10568
rect 4618 10240 4674 10296
rect 4904 10906 4960 10908
rect 4984 10906 5040 10908
rect 5064 10906 5120 10908
rect 5144 10906 5200 10908
rect 4904 10854 4950 10906
rect 4950 10854 4960 10906
rect 4984 10854 5014 10906
rect 5014 10854 5026 10906
rect 5026 10854 5040 10906
rect 5064 10854 5078 10906
rect 5078 10854 5090 10906
rect 5090 10854 5120 10906
rect 5144 10854 5154 10906
rect 5154 10854 5200 10906
rect 4904 10852 4960 10854
rect 4984 10852 5040 10854
rect 5064 10852 5120 10854
rect 5144 10852 5200 10854
rect 4894 10512 4950 10568
rect 4904 9818 4960 9820
rect 4984 9818 5040 9820
rect 5064 9818 5120 9820
rect 5144 9818 5200 9820
rect 4904 9766 4950 9818
rect 4950 9766 4960 9818
rect 4984 9766 5014 9818
rect 5014 9766 5026 9818
rect 5026 9766 5040 9818
rect 5064 9766 5078 9818
rect 5078 9766 5090 9818
rect 5090 9766 5120 9818
rect 5144 9766 5154 9818
rect 5154 9766 5200 9818
rect 4904 9764 4960 9766
rect 4984 9764 5040 9766
rect 5064 9764 5120 9766
rect 5144 9764 5200 9766
rect 4904 8730 4960 8732
rect 4984 8730 5040 8732
rect 5064 8730 5120 8732
rect 5144 8730 5200 8732
rect 4904 8678 4950 8730
rect 4950 8678 4960 8730
rect 4984 8678 5014 8730
rect 5014 8678 5026 8730
rect 5026 8678 5040 8730
rect 5064 8678 5078 8730
rect 5078 8678 5090 8730
rect 5090 8678 5120 8730
rect 5144 8678 5154 8730
rect 5154 8678 5200 8730
rect 4904 8676 4960 8678
rect 4984 8676 5040 8678
rect 5064 8676 5120 8678
rect 5144 8676 5200 8678
rect 5446 19760 5502 19816
rect 5630 19624 5686 19680
rect 5814 20168 5870 20204
rect 6090 19896 6146 19952
rect 5906 19488 5962 19544
rect 5722 18808 5778 18864
rect 5630 18128 5686 18184
rect 5446 16768 5502 16824
rect 5354 14456 5410 14512
rect 5630 13640 5686 13696
rect 5446 12688 5502 12744
rect 6090 18944 6146 19000
rect 5814 13368 5870 13424
rect 5814 13096 5870 13152
rect 6642 19760 6698 19816
rect 6550 19352 6606 19408
rect 6274 18264 6330 18320
rect 6366 17856 6422 17912
rect 6550 17992 6606 18048
rect 6366 17448 6422 17504
rect 6458 17176 6514 17232
rect 6090 15136 6146 15192
rect 5446 8608 5502 8664
rect 5078 8356 5134 8392
rect 5078 8336 5080 8356
rect 5080 8336 5132 8356
rect 5132 8336 5134 8356
rect 4802 7812 4858 7848
rect 4802 7792 4804 7812
rect 4804 7792 4856 7812
rect 4856 7792 4858 7812
rect 4904 7642 4960 7644
rect 4984 7642 5040 7644
rect 5064 7642 5120 7644
rect 5144 7642 5200 7644
rect 4904 7590 4950 7642
rect 4950 7590 4960 7642
rect 4984 7590 5014 7642
rect 5014 7590 5026 7642
rect 5026 7590 5040 7642
rect 5064 7590 5078 7642
rect 5078 7590 5090 7642
rect 5090 7590 5120 7642
rect 5144 7590 5154 7642
rect 5154 7590 5200 7642
rect 4904 7588 4960 7590
rect 4984 7588 5040 7590
rect 5064 7588 5120 7590
rect 5144 7588 5200 7590
rect 4904 6554 4960 6556
rect 4984 6554 5040 6556
rect 5064 6554 5120 6556
rect 5144 6554 5200 6556
rect 4904 6502 4950 6554
rect 4950 6502 4960 6554
rect 4984 6502 5014 6554
rect 5014 6502 5026 6554
rect 5026 6502 5040 6554
rect 5064 6502 5078 6554
rect 5078 6502 5090 6554
rect 5090 6502 5120 6554
rect 5144 6502 5154 6554
rect 5154 6502 5200 6554
rect 4904 6500 4960 6502
rect 4984 6500 5040 6502
rect 5064 6500 5120 6502
rect 5144 6500 5200 6502
rect 4904 5466 4960 5468
rect 4984 5466 5040 5468
rect 5064 5466 5120 5468
rect 5144 5466 5200 5468
rect 4904 5414 4950 5466
rect 4950 5414 4960 5466
rect 4984 5414 5014 5466
rect 5014 5414 5026 5466
rect 5026 5414 5040 5466
rect 5064 5414 5078 5466
rect 5078 5414 5090 5466
rect 5090 5414 5120 5466
rect 5144 5414 5154 5466
rect 5154 5414 5200 5466
rect 4904 5412 4960 5414
rect 4984 5412 5040 5414
rect 5064 5412 5120 5414
rect 5144 5412 5200 5414
rect 5170 5072 5226 5128
rect 4904 4378 4960 4380
rect 4984 4378 5040 4380
rect 5064 4378 5120 4380
rect 5144 4378 5200 4380
rect 4904 4326 4950 4378
rect 4950 4326 4960 4378
rect 4984 4326 5014 4378
rect 5014 4326 5026 4378
rect 5026 4326 5040 4378
rect 5064 4326 5078 4378
rect 5078 4326 5090 4378
rect 5090 4326 5120 4378
rect 5144 4326 5154 4378
rect 5154 4326 5200 4378
rect 4904 4324 4960 4326
rect 4984 4324 5040 4326
rect 5064 4324 5120 4326
rect 5144 4324 5200 4326
rect 4802 3984 4858 4040
rect 4434 2760 4490 2816
rect 4904 3290 4960 3292
rect 4984 3290 5040 3292
rect 5064 3290 5120 3292
rect 5144 3290 5200 3292
rect 4904 3238 4950 3290
rect 4950 3238 4960 3290
rect 4984 3238 5014 3290
rect 5014 3238 5026 3290
rect 5026 3238 5040 3290
rect 5064 3238 5078 3290
rect 5078 3238 5090 3290
rect 5090 3238 5120 3290
rect 5144 3238 5154 3290
rect 5154 3238 5200 3290
rect 4904 3236 4960 3238
rect 4984 3236 5040 3238
rect 5064 3236 5120 3238
rect 5144 3236 5200 3238
rect 4904 2202 4960 2204
rect 4984 2202 5040 2204
rect 5064 2202 5120 2204
rect 5144 2202 5200 2204
rect 4904 2150 4950 2202
rect 4950 2150 4960 2202
rect 4984 2150 5014 2202
rect 5014 2150 5026 2202
rect 5026 2150 5040 2202
rect 5064 2150 5078 2202
rect 5078 2150 5090 2202
rect 5090 2150 5120 2202
rect 5144 2150 5154 2202
rect 5154 2150 5200 2202
rect 4904 2148 4960 2150
rect 4984 2148 5040 2150
rect 5064 2148 5120 2150
rect 5144 2148 5200 2150
rect 5170 1808 5226 1864
rect 4904 1114 4960 1116
rect 4984 1114 5040 1116
rect 5064 1114 5120 1116
rect 5144 1114 5200 1116
rect 4904 1062 4950 1114
rect 4950 1062 4960 1114
rect 4984 1062 5014 1114
rect 5014 1062 5026 1114
rect 5026 1062 5040 1114
rect 5064 1062 5078 1114
rect 5078 1062 5090 1114
rect 5090 1062 5120 1114
rect 5144 1062 5154 1114
rect 5154 1062 5200 1114
rect 4904 1060 4960 1062
rect 4984 1060 5040 1062
rect 5064 1060 5120 1062
rect 5144 1060 5200 1062
rect 5722 9968 5778 10024
rect 5630 7384 5686 7440
rect 5538 6024 5594 6080
rect 5538 5480 5594 5536
rect 5538 4528 5594 4584
rect 5446 3168 5502 3224
rect 5998 11872 6054 11928
rect 5998 10240 6054 10296
rect 5998 10104 6054 10160
rect 6274 15544 6330 15600
rect 6182 14592 6238 14648
rect 6182 12960 6238 13016
rect 6182 12280 6238 12336
rect 6878 21242 6934 21244
rect 6958 21242 7014 21244
rect 7038 21242 7094 21244
rect 7118 21242 7174 21244
rect 6878 21190 6924 21242
rect 6924 21190 6934 21242
rect 6958 21190 6988 21242
rect 6988 21190 7000 21242
rect 7000 21190 7014 21242
rect 7038 21190 7052 21242
rect 7052 21190 7064 21242
rect 7064 21190 7094 21242
rect 7118 21190 7128 21242
rect 7128 21190 7174 21242
rect 6878 21188 6934 21190
rect 6958 21188 7014 21190
rect 7038 21188 7094 21190
rect 7118 21188 7174 21190
rect 6878 20154 6934 20156
rect 6958 20154 7014 20156
rect 7038 20154 7094 20156
rect 7118 20154 7174 20156
rect 6878 20102 6924 20154
rect 6924 20102 6934 20154
rect 6958 20102 6988 20154
rect 6988 20102 7000 20154
rect 7000 20102 7014 20154
rect 7038 20102 7052 20154
rect 7052 20102 7064 20154
rect 7064 20102 7094 20154
rect 7118 20102 7128 20154
rect 7128 20102 7174 20154
rect 6878 20100 6934 20102
rect 6958 20100 7014 20102
rect 7038 20100 7094 20102
rect 7118 20100 7174 20102
rect 6878 19066 6934 19068
rect 6958 19066 7014 19068
rect 7038 19066 7094 19068
rect 7118 19066 7174 19068
rect 6878 19014 6924 19066
rect 6924 19014 6934 19066
rect 6958 19014 6988 19066
rect 6988 19014 7000 19066
rect 7000 19014 7014 19066
rect 7038 19014 7052 19066
rect 7052 19014 7064 19066
rect 7064 19014 7094 19066
rect 7118 19014 7128 19066
rect 7128 19014 7174 19066
rect 6878 19012 6934 19014
rect 6958 19012 7014 19014
rect 7038 19012 7094 19014
rect 7118 19012 7174 19014
rect 7654 18536 7710 18592
rect 7102 18264 7158 18320
rect 6878 17978 6934 17980
rect 6958 17978 7014 17980
rect 7038 17978 7094 17980
rect 7118 17978 7174 17980
rect 6878 17926 6924 17978
rect 6924 17926 6934 17978
rect 6958 17926 6988 17978
rect 6988 17926 7000 17978
rect 7000 17926 7014 17978
rect 7038 17926 7052 17978
rect 7052 17926 7064 17978
rect 7064 17926 7094 17978
rect 7118 17926 7128 17978
rect 7128 17926 7174 17978
rect 6878 17924 6934 17926
rect 6958 17924 7014 17926
rect 7038 17924 7094 17926
rect 7118 17924 7174 17926
rect 7102 17604 7158 17640
rect 7102 17584 7104 17604
rect 7104 17584 7156 17604
rect 7156 17584 7158 17604
rect 6878 16890 6934 16892
rect 6958 16890 7014 16892
rect 7038 16890 7094 16892
rect 7118 16890 7174 16892
rect 6878 16838 6924 16890
rect 6924 16838 6934 16890
rect 6958 16838 6988 16890
rect 6988 16838 7000 16890
rect 7000 16838 7014 16890
rect 7038 16838 7052 16890
rect 7052 16838 7064 16890
rect 7064 16838 7094 16890
rect 7118 16838 7128 16890
rect 7128 16838 7174 16890
rect 6878 16836 6934 16838
rect 6958 16836 7014 16838
rect 7038 16836 7094 16838
rect 7118 16836 7174 16838
rect 6918 16632 6974 16688
rect 6734 16360 6790 16416
rect 6642 16224 6698 16280
rect 6642 15272 6698 15328
rect 6458 14864 6514 14920
rect 7654 17448 7710 17504
rect 7378 17312 7434 17368
rect 7470 16768 7526 16824
rect 7378 16496 7434 16552
rect 7286 16224 7342 16280
rect 6878 15802 6934 15804
rect 6958 15802 7014 15804
rect 7038 15802 7094 15804
rect 7118 15802 7174 15804
rect 6878 15750 6924 15802
rect 6924 15750 6934 15802
rect 6958 15750 6988 15802
rect 6988 15750 7000 15802
rect 7000 15750 7014 15802
rect 7038 15750 7052 15802
rect 7052 15750 7064 15802
rect 7064 15750 7094 15802
rect 7118 15750 7128 15802
rect 7128 15750 7174 15802
rect 6878 15748 6934 15750
rect 6958 15748 7014 15750
rect 7038 15748 7094 15750
rect 7118 15748 7174 15750
rect 7194 15020 7250 15056
rect 7194 15000 7196 15020
rect 7196 15000 7248 15020
rect 7248 15000 7250 15020
rect 6878 14714 6934 14716
rect 6958 14714 7014 14716
rect 7038 14714 7094 14716
rect 7118 14714 7174 14716
rect 6878 14662 6924 14714
rect 6924 14662 6934 14714
rect 6958 14662 6988 14714
rect 6988 14662 7000 14714
rect 7000 14662 7014 14714
rect 7038 14662 7052 14714
rect 7052 14662 7064 14714
rect 7064 14662 7094 14714
rect 7118 14662 7128 14714
rect 7128 14662 7174 14714
rect 6878 14660 6934 14662
rect 6958 14660 7014 14662
rect 7038 14660 7094 14662
rect 7118 14660 7174 14662
rect 6734 14592 6790 14648
rect 6458 14456 6514 14512
rect 6366 13232 6422 13288
rect 6366 12824 6422 12880
rect 6366 12708 6422 12744
rect 6366 12688 6368 12708
rect 6368 12688 6420 12708
rect 6420 12688 6422 12708
rect 6182 10376 6238 10432
rect 6090 9288 6146 9344
rect 6734 14184 6790 14240
rect 7470 15000 7526 15056
rect 6878 13626 6934 13628
rect 6958 13626 7014 13628
rect 7038 13626 7094 13628
rect 7118 13626 7174 13628
rect 6878 13574 6924 13626
rect 6924 13574 6934 13626
rect 6958 13574 6988 13626
rect 6988 13574 7000 13626
rect 7000 13574 7014 13626
rect 7038 13574 7052 13626
rect 7052 13574 7064 13626
rect 7064 13574 7094 13626
rect 7118 13574 7128 13626
rect 7128 13574 7174 13626
rect 6878 13572 6934 13574
rect 6958 13572 7014 13574
rect 7038 13572 7094 13574
rect 7118 13572 7174 13574
rect 6642 13096 6698 13152
rect 6458 12280 6514 12336
rect 6182 9016 6238 9072
rect 5814 4392 5870 4448
rect 5814 3712 5870 3768
rect 6274 8880 6330 8936
rect 6182 7928 6238 7984
rect 6182 7520 6238 7576
rect 6274 6568 6330 6624
rect 5998 3440 6054 3496
rect 5998 3032 6054 3088
rect 5998 2216 6054 2272
rect 6182 3032 6238 3088
rect 6090 2080 6146 2136
rect 7010 12960 7066 13016
rect 7010 12688 7066 12744
rect 7470 14456 7526 14512
rect 7378 12824 7434 12880
rect 7562 12860 7564 12880
rect 7564 12860 7616 12880
rect 7616 12860 7618 12880
rect 7562 12824 7618 12860
rect 6878 12538 6934 12540
rect 6958 12538 7014 12540
rect 7038 12538 7094 12540
rect 7118 12538 7174 12540
rect 6878 12486 6924 12538
rect 6924 12486 6934 12538
rect 6958 12486 6988 12538
rect 6988 12486 7000 12538
rect 7000 12486 7014 12538
rect 7038 12486 7052 12538
rect 7052 12486 7064 12538
rect 7064 12486 7094 12538
rect 7118 12486 7128 12538
rect 7128 12486 7174 12538
rect 6878 12484 6934 12486
rect 6958 12484 7014 12486
rect 7038 12484 7094 12486
rect 7118 12484 7174 12486
rect 6734 12144 6790 12200
rect 6918 12180 6920 12200
rect 6920 12180 6972 12200
rect 6972 12180 6974 12200
rect 6918 12144 6974 12180
rect 6642 11736 6698 11792
rect 6878 11450 6934 11452
rect 6958 11450 7014 11452
rect 7038 11450 7094 11452
rect 7118 11450 7174 11452
rect 6878 11398 6924 11450
rect 6924 11398 6934 11450
rect 6958 11398 6988 11450
rect 6988 11398 7000 11450
rect 7000 11398 7014 11450
rect 7038 11398 7052 11450
rect 7052 11398 7064 11450
rect 7064 11398 7094 11450
rect 7118 11398 7128 11450
rect 7128 11398 7174 11450
rect 6878 11396 6934 11398
rect 6958 11396 7014 11398
rect 7038 11396 7094 11398
rect 7118 11396 7174 11398
rect 7102 11192 7158 11248
rect 6878 10362 6934 10364
rect 6958 10362 7014 10364
rect 7038 10362 7094 10364
rect 7118 10362 7174 10364
rect 6878 10310 6924 10362
rect 6924 10310 6934 10362
rect 6958 10310 6988 10362
rect 6988 10310 7000 10362
rect 7000 10310 7014 10362
rect 7038 10310 7052 10362
rect 7052 10310 7064 10362
rect 7064 10310 7094 10362
rect 7118 10310 7128 10362
rect 7128 10310 7174 10362
rect 6878 10308 6934 10310
rect 6958 10308 7014 10310
rect 7038 10308 7094 10310
rect 7118 10308 7174 10310
rect 7470 12552 7526 12608
rect 7562 12280 7618 12336
rect 7378 11328 7434 11384
rect 6826 9696 6882 9752
rect 6878 9274 6934 9276
rect 6958 9274 7014 9276
rect 7038 9274 7094 9276
rect 7118 9274 7174 9276
rect 6878 9222 6924 9274
rect 6924 9222 6934 9274
rect 6958 9222 6988 9274
rect 6988 9222 7000 9274
rect 7000 9222 7014 9274
rect 7038 9222 7052 9274
rect 7052 9222 7064 9274
rect 7064 9222 7094 9274
rect 7118 9222 7128 9274
rect 7128 9222 7174 9274
rect 6878 9220 6934 9222
rect 6958 9220 7014 9222
rect 7038 9220 7094 9222
rect 7118 9220 7174 9222
rect 6734 8744 6790 8800
rect 6550 7928 6606 7984
rect 6878 8186 6934 8188
rect 6958 8186 7014 8188
rect 7038 8186 7094 8188
rect 7118 8186 7174 8188
rect 6878 8134 6924 8186
rect 6924 8134 6934 8186
rect 6958 8134 6988 8186
rect 6988 8134 7000 8186
rect 7000 8134 7014 8186
rect 7038 8134 7052 8186
rect 7052 8134 7064 8186
rect 7064 8134 7094 8186
rect 7118 8134 7128 8186
rect 7128 8134 7174 8186
rect 6878 8132 6934 8134
rect 6958 8132 7014 8134
rect 7038 8132 7094 8134
rect 7118 8132 7174 8134
rect 7010 7404 7066 7440
rect 7010 7384 7012 7404
rect 7012 7384 7064 7404
rect 7064 7384 7066 7404
rect 6878 7098 6934 7100
rect 6958 7098 7014 7100
rect 7038 7098 7094 7100
rect 7118 7098 7174 7100
rect 6878 7046 6924 7098
rect 6924 7046 6934 7098
rect 6958 7046 6988 7098
rect 6988 7046 7000 7098
rect 7000 7046 7014 7098
rect 7038 7046 7052 7098
rect 7052 7046 7064 7098
rect 7064 7046 7094 7098
rect 7118 7046 7128 7098
rect 7128 7046 7174 7098
rect 6878 7044 6934 7046
rect 6958 7044 7014 7046
rect 7038 7044 7094 7046
rect 7118 7044 7174 7046
rect 7194 6432 7250 6488
rect 7102 6316 7158 6352
rect 7102 6296 7104 6316
rect 7104 6296 7156 6316
rect 7156 6296 7158 6316
rect 6878 6010 6934 6012
rect 6958 6010 7014 6012
rect 7038 6010 7094 6012
rect 7118 6010 7174 6012
rect 6878 5958 6924 6010
rect 6924 5958 6934 6010
rect 6958 5958 6988 6010
rect 6988 5958 7000 6010
rect 7000 5958 7014 6010
rect 7038 5958 7052 6010
rect 7052 5958 7064 6010
rect 7064 5958 7094 6010
rect 7118 5958 7128 6010
rect 7128 5958 7174 6010
rect 6878 5956 6934 5958
rect 6958 5956 7014 5958
rect 7038 5956 7094 5958
rect 7118 5956 7174 5958
rect 6458 5364 6514 5400
rect 6458 5344 6460 5364
rect 6460 5344 6512 5364
rect 6512 5344 6514 5364
rect 6734 5344 6790 5400
rect 7010 5344 7066 5400
rect 6642 5108 6644 5128
rect 6644 5108 6696 5128
rect 6696 5108 6698 5128
rect 6642 5072 6698 5108
rect 6642 4664 6698 4720
rect 6458 3848 6514 3904
rect 6878 4922 6934 4924
rect 6958 4922 7014 4924
rect 7038 4922 7094 4924
rect 7118 4922 7174 4924
rect 6878 4870 6924 4922
rect 6924 4870 6934 4922
rect 6958 4870 6988 4922
rect 6988 4870 7000 4922
rect 7000 4870 7014 4922
rect 7038 4870 7052 4922
rect 7052 4870 7064 4922
rect 7064 4870 7094 4922
rect 7118 4870 7128 4922
rect 7128 4870 7174 4922
rect 6878 4868 6934 4870
rect 6958 4868 7014 4870
rect 7038 4868 7094 4870
rect 7118 4868 7174 4870
rect 6918 4664 6974 4720
rect 6826 4528 6882 4584
rect 6642 3884 6644 3904
rect 6644 3884 6696 3904
rect 6696 3884 6698 3904
rect 6642 3848 6698 3884
rect 6878 3834 6934 3836
rect 6958 3834 7014 3836
rect 7038 3834 7094 3836
rect 7118 3834 7174 3836
rect 6878 3782 6924 3834
rect 6924 3782 6934 3834
rect 6958 3782 6988 3834
rect 6988 3782 7000 3834
rect 7000 3782 7014 3834
rect 7038 3782 7052 3834
rect 7052 3782 7064 3834
rect 7064 3782 7094 3834
rect 7118 3782 7128 3834
rect 7128 3782 7174 3834
rect 6878 3780 6934 3782
rect 6958 3780 7014 3782
rect 7038 3780 7094 3782
rect 7118 3780 7174 3782
rect 6550 3168 6606 3224
rect 6274 1536 6330 1592
rect 6182 856 6238 912
rect 7010 3304 7066 3360
rect 7378 6024 7434 6080
rect 7378 4392 7434 4448
rect 7378 3848 7434 3904
rect 7562 6432 7618 6488
rect 7930 18264 7986 18320
rect 8482 18844 8484 18864
rect 8484 18844 8536 18864
rect 8536 18844 8538 18864
rect 8482 18808 8538 18844
rect 8482 18672 8538 18728
rect 8852 21786 8908 21788
rect 8932 21786 8988 21788
rect 9012 21786 9068 21788
rect 9092 21786 9148 21788
rect 8852 21734 8898 21786
rect 8898 21734 8908 21786
rect 8932 21734 8962 21786
rect 8962 21734 8974 21786
rect 8974 21734 8988 21786
rect 9012 21734 9026 21786
rect 9026 21734 9038 21786
rect 9038 21734 9068 21786
rect 9092 21734 9102 21786
rect 9102 21734 9148 21786
rect 8852 21732 8908 21734
rect 8932 21732 8988 21734
rect 9012 21732 9068 21734
rect 9092 21732 9148 21734
rect 12800 21786 12856 21788
rect 12880 21786 12936 21788
rect 12960 21786 13016 21788
rect 13040 21786 13096 21788
rect 12800 21734 12846 21786
rect 12846 21734 12856 21786
rect 12880 21734 12910 21786
rect 12910 21734 12922 21786
rect 12922 21734 12936 21786
rect 12960 21734 12974 21786
rect 12974 21734 12986 21786
rect 12986 21734 13016 21786
rect 13040 21734 13050 21786
rect 13050 21734 13096 21786
rect 12800 21732 12856 21734
rect 12880 21732 12936 21734
rect 12960 21732 13016 21734
rect 13040 21732 13096 21734
rect 8852 20698 8908 20700
rect 8932 20698 8988 20700
rect 9012 20698 9068 20700
rect 9092 20698 9148 20700
rect 8852 20646 8898 20698
rect 8898 20646 8908 20698
rect 8932 20646 8962 20698
rect 8962 20646 8974 20698
rect 8974 20646 8988 20698
rect 9012 20646 9026 20698
rect 9026 20646 9038 20698
rect 9038 20646 9068 20698
rect 9092 20646 9102 20698
rect 9102 20646 9148 20698
rect 8852 20644 8908 20646
rect 8932 20644 8988 20646
rect 9012 20644 9068 20646
rect 9092 20644 9148 20646
rect 8666 19624 8722 19680
rect 7930 17856 7986 17912
rect 8114 18028 8116 18048
rect 8116 18028 8168 18048
rect 8168 18028 8170 18048
rect 8114 17992 8170 18028
rect 8206 17448 8262 17504
rect 7930 16768 7986 16824
rect 7838 16632 7894 16688
rect 8022 16244 8078 16280
rect 8022 16224 8024 16244
rect 8024 16224 8076 16244
rect 8076 16224 8078 16244
rect 8298 17312 8354 17368
rect 8298 16532 8300 16552
rect 8300 16532 8352 16552
rect 8352 16532 8354 16552
rect 8298 16496 8354 16532
rect 7746 15816 7802 15872
rect 7746 13776 7802 13832
rect 7746 12960 7802 13016
rect 7746 12688 7802 12744
rect 7930 12688 7986 12744
rect 8022 12552 8078 12608
rect 8206 13504 8262 13560
rect 7930 9696 7986 9752
rect 8206 12144 8262 12200
rect 8206 11328 8262 11384
rect 8114 9968 8170 10024
rect 7930 7420 7932 7440
rect 7932 7420 7984 7440
rect 7984 7420 7986 7440
rect 7930 7384 7986 7420
rect 8022 7112 8078 7168
rect 8114 6704 8170 6760
rect 8574 17448 8630 17504
rect 8482 16904 8538 16960
rect 8852 19610 8908 19612
rect 8932 19610 8988 19612
rect 9012 19610 9068 19612
rect 9092 19610 9148 19612
rect 8852 19558 8898 19610
rect 8898 19558 8908 19610
rect 8932 19558 8962 19610
rect 8962 19558 8974 19610
rect 8974 19558 8988 19610
rect 9012 19558 9026 19610
rect 9026 19558 9038 19610
rect 9038 19558 9068 19610
rect 9092 19558 9102 19610
rect 9102 19558 9148 19610
rect 8852 19556 8908 19558
rect 8932 19556 8988 19558
rect 9012 19556 9068 19558
rect 9092 19556 9148 19558
rect 9218 19352 9274 19408
rect 8852 18522 8908 18524
rect 8932 18522 8988 18524
rect 9012 18522 9068 18524
rect 9092 18522 9148 18524
rect 8852 18470 8898 18522
rect 8898 18470 8908 18522
rect 8932 18470 8962 18522
rect 8962 18470 8974 18522
rect 8974 18470 8988 18522
rect 9012 18470 9026 18522
rect 9026 18470 9038 18522
rect 9038 18470 9068 18522
rect 9092 18470 9102 18522
rect 9102 18470 9148 18522
rect 8852 18468 8908 18470
rect 8932 18468 8988 18470
rect 9012 18468 9068 18470
rect 9092 18468 9148 18470
rect 8482 16224 8538 16280
rect 8482 14864 8538 14920
rect 10826 21242 10882 21244
rect 10906 21242 10962 21244
rect 10986 21242 11042 21244
rect 11066 21242 11122 21244
rect 10826 21190 10872 21242
rect 10872 21190 10882 21242
rect 10906 21190 10936 21242
rect 10936 21190 10948 21242
rect 10948 21190 10962 21242
rect 10986 21190 11000 21242
rect 11000 21190 11012 21242
rect 11012 21190 11042 21242
rect 11066 21190 11076 21242
rect 11076 21190 11122 21242
rect 10826 21188 10882 21190
rect 10906 21188 10962 21190
rect 10986 21188 11042 21190
rect 11066 21188 11122 21190
rect 9494 18264 9550 18320
rect 9678 17992 9734 18048
rect 9402 17720 9458 17776
rect 8852 17434 8908 17436
rect 8932 17434 8988 17436
rect 9012 17434 9068 17436
rect 9092 17434 9148 17436
rect 8852 17382 8898 17434
rect 8898 17382 8908 17434
rect 8932 17382 8962 17434
rect 8962 17382 8974 17434
rect 8974 17382 8988 17434
rect 9012 17382 9026 17434
rect 9026 17382 9038 17434
rect 9038 17382 9068 17434
rect 9092 17382 9102 17434
rect 9102 17382 9148 17434
rect 8852 17380 8908 17382
rect 8932 17380 8988 17382
rect 9012 17380 9068 17382
rect 9092 17380 9148 17382
rect 9034 17040 9090 17096
rect 8852 16346 8908 16348
rect 8932 16346 8988 16348
rect 9012 16346 9068 16348
rect 9092 16346 9148 16348
rect 8852 16294 8898 16346
rect 8898 16294 8908 16346
rect 8932 16294 8962 16346
rect 8962 16294 8974 16346
rect 8974 16294 8988 16346
rect 9012 16294 9026 16346
rect 9026 16294 9038 16346
rect 9038 16294 9068 16346
rect 9092 16294 9102 16346
rect 9102 16294 9148 16346
rect 8852 16292 8908 16294
rect 8932 16292 8988 16294
rect 9012 16292 9068 16294
rect 9092 16292 9148 16294
rect 9034 15816 9090 15872
rect 8942 15408 8998 15464
rect 9678 17040 9734 17096
rect 9862 17448 9918 17504
rect 9494 16904 9550 16960
rect 9678 16940 9680 16960
rect 9680 16940 9732 16960
rect 9732 16940 9734 16960
rect 9678 16904 9734 16940
rect 9310 16224 9366 16280
rect 9310 15816 9366 15872
rect 9678 16396 9680 16416
rect 9680 16396 9732 16416
rect 9732 16396 9734 16416
rect 9678 16360 9734 16396
rect 10046 17312 10102 17368
rect 10046 17040 10102 17096
rect 9954 16360 10010 16416
rect 9770 16088 9826 16144
rect 9218 15408 9274 15464
rect 8852 15258 8908 15260
rect 8932 15258 8988 15260
rect 9012 15258 9068 15260
rect 9092 15258 9148 15260
rect 8852 15206 8898 15258
rect 8898 15206 8908 15258
rect 8932 15206 8962 15258
rect 8962 15206 8974 15258
rect 8974 15206 8988 15258
rect 9012 15206 9026 15258
rect 9026 15206 9038 15258
rect 9038 15206 9068 15258
rect 9092 15206 9102 15258
rect 9102 15206 9148 15258
rect 8852 15204 8908 15206
rect 8932 15204 8988 15206
rect 9012 15204 9068 15206
rect 9092 15204 9148 15206
rect 8758 14492 8760 14512
rect 8760 14492 8812 14512
rect 8812 14492 8814 14512
rect 8758 14456 8814 14492
rect 9126 14728 9182 14784
rect 9310 14864 9366 14920
rect 9126 14492 9128 14512
rect 9128 14492 9180 14512
rect 9180 14492 9182 14512
rect 9126 14456 9182 14492
rect 8574 14184 8630 14240
rect 8482 12960 8538 13016
rect 8852 14170 8908 14172
rect 8932 14170 8988 14172
rect 9012 14170 9068 14172
rect 9092 14170 9148 14172
rect 8852 14118 8898 14170
rect 8898 14118 8908 14170
rect 8932 14118 8962 14170
rect 8962 14118 8974 14170
rect 8974 14118 8988 14170
rect 9012 14118 9026 14170
rect 9026 14118 9038 14170
rect 9038 14118 9068 14170
rect 9092 14118 9102 14170
rect 9102 14118 9148 14170
rect 8852 14116 8908 14118
rect 8932 14116 8988 14118
rect 9012 14116 9068 14118
rect 9092 14116 9148 14118
rect 8850 13776 8906 13832
rect 8942 13640 8998 13696
rect 9126 13504 9182 13560
rect 8666 12960 8722 13016
rect 8574 12144 8630 12200
rect 8482 10920 8538 10976
rect 8390 10648 8446 10704
rect 8298 10240 8354 10296
rect 8298 8336 8354 8392
rect 8206 6432 8262 6488
rect 6642 2488 6698 2544
rect 7286 2760 7342 2816
rect 6878 2746 6934 2748
rect 6958 2746 7014 2748
rect 7038 2746 7094 2748
rect 7118 2746 7174 2748
rect 6878 2694 6924 2746
rect 6924 2694 6934 2746
rect 6958 2694 6988 2746
rect 6988 2694 7000 2746
rect 7000 2694 7014 2746
rect 7038 2694 7052 2746
rect 7052 2694 7064 2746
rect 7064 2694 7094 2746
rect 7118 2694 7128 2746
rect 7128 2694 7174 2746
rect 6878 2692 6934 2694
rect 6958 2692 7014 2694
rect 7038 2692 7094 2694
rect 7118 2692 7174 2694
rect 7562 2624 7618 2680
rect 7654 2352 7710 2408
rect 6878 1658 6934 1660
rect 6958 1658 7014 1660
rect 7038 1658 7094 1660
rect 7118 1658 7174 1660
rect 6878 1606 6924 1658
rect 6924 1606 6934 1658
rect 6958 1606 6988 1658
rect 6988 1606 7000 1658
rect 7000 1606 7014 1658
rect 7038 1606 7052 1658
rect 7052 1606 7064 1658
rect 7064 1606 7094 1658
rect 7118 1606 7128 1658
rect 7128 1606 7174 1658
rect 6878 1604 6934 1606
rect 6958 1604 7014 1606
rect 7038 1604 7094 1606
rect 7118 1604 7174 1606
rect 7286 1536 7342 1592
rect 6826 1400 6882 1456
rect 7010 1400 7066 1456
rect 6458 1128 6514 1184
rect 7838 1672 7894 1728
rect 8022 5072 8078 5128
rect 8022 4256 8078 4312
rect 8022 3712 8078 3768
rect 8298 5480 8354 5536
rect 8298 4528 8354 4584
rect 8022 3440 8078 3496
rect 8206 3304 8262 3360
rect 8852 13082 8908 13084
rect 8932 13082 8988 13084
rect 9012 13082 9068 13084
rect 9092 13082 9148 13084
rect 8852 13030 8898 13082
rect 8898 13030 8908 13082
rect 8932 13030 8962 13082
rect 8962 13030 8974 13082
rect 8974 13030 8988 13082
rect 9012 13030 9026 13082
rect 9026 13030 9038 13082
rect 9038 13030 9068 13082
rect 9092 13030 9102 13082
rect 9102 13030 9148 13082
rect 8852 13028 8908 13030
rect 8932 13028 8988 13030
rect 9012 13028 9068 13030
rect 9092 13028 9148 13030
rect 9126 12688 9182 12744
rect 9034 12144 9090 12200
rect 9494 15408 9550 15464
rect 9402 14220 9404 14240
rect 9404 14220 9456 14240
rect 9456 14220 9458 14240
rect 9402 14184 9458 14220
rect 9218 12416 9274 12472
rect 8852 11994 8908 11996
rect 8932 11994 8988 11996
rect 9012 11994 9068 11996
rect 9092 11994 9148 11996
rect 8852 11942 8898 11994
rect 8898 11942 8908 11994
rect 8932 11942 8962 11994
rect 8962 11942 8974 11994
rect 8974 11942 8988 11994
rect 9012 11942 9026 11994
rect 9026 11942 9038 11994
rect 9038 11942 9068 11994
rect 9092 11942 9102 11994
rect 9102 11942 9148 11994
rect 8852 11940 8908 11942
rect 8932 11940 8988 11942
rect 9012 11940 9068 11942
rect 9092 11940 9148 11942
rect 9034 11076 9090 11112
rect 9034 11056 9036 11076
rect 9036 11056 9088 11076
rect 9088 11056 9090 11076
rect 8852 10906 8908 10908
rect 8932 10906 8988 10908
rect 9012 10906 9068 10908
rect 9092 10906 9148 10908
rect 8852 10854 8898 10906
rect 8898 10854 8908 10906
rect 8932 10854 8962 10906
rect 8962 10854 8974 10906
rect 8974 10854 8988 10906
rect 9012 10854 9026 10906
rect 9026 10854 9038 10906
rect 9038 10854 9068 10906
rect 9092 10854 9102 10906
rect 9102 10854 9148 10906
rect 8852 10852 8908 10854
rect 8932 10852 8988 10854
rect 9012 10852 9068 10854
rect 9092 10852 9148 10854
rect 9034 10648 9090 10704
rect 9494 13096 9550 13152
rect 9954 15000 10010 15056
rect 9862 13676 9864 13696
rect 9864 13676 9916 13696
rect 9916 13676 9918 13696
rect 9862 13640 9918 13676
rect 9954 12960 10010 13016
rect 9770 12688 9826 12744
rect 9586 12280 9642 12336
rect 9770 12280 9826 12336
rect 9402 12008 9458 12064
rect 9586 12144 9642 12200
rect 9586 12008 9642 12064
rect 9310 11192 9366 11248
rect 8574 9868 8576 9888
rect 8576 9868 8628 9888
rect 8628 9868 8630 9888
rect 8574 9832 8630 9868
rect 9218 9968 9274 10024
rect 8852 9818 8908 9820
rect 8932 9818 8988 9820
rect 9012 9818 9068 9820
rect 9092 9818 9148 9820
rect 8852 9766 8898 9818
rect 8898 9766 8908 9818
rect 8932 9766 8962 9818
rect 8962 9766 8974 9818
rect 8974 9766 8988 9818
rect 9012 9766 9026 9818
rect 9026 9766 9038 9818
rect 9038 9766 9068 9818
rect 9092 9766 9102 9818
rect 9102 9766 9148 9818
rect 8852 9764 8908 9766
rect 8932 9764 8988 9766
rect 9012 9764 9068 9766
rect 9092 9764 9148 9766
rect 8758 9016 8814 9072
rect 8666 8744 8722 8800
rect 8852 8730 8908 8732
rect 8932 8730 8988 8732
rect 9012 8730 9068 8732
rect 9092 8730 9148 8732
rect 8852 8678 8898 8730
rect 8898 8678 8908 8730
rect 8932 8678 8962 8730
rect 8962 8678 8974 8730
rect 8974 8678 8988 8730
rect 9012 8678 9026 8730
rect 9026 8678 9038 8730
rect 9038 8678 9068 8730
rect 9092 8678 9102 8730
rect 9102 8678 9148 8730
rect 8852 8676 8908 8678
rect 8932 8676 8988 8678
rect 9012 8676 9068 8678
rect 9092 8676 9148 8678
rect 8666 8608 8722 8664
rect 8758 8200 8814 8256
rect 9034 8200 9090 8256
rect 8574 7656 8630 7712
rect 8482 5344 8538 5400
rect 8482 3440 8538 3496
rect 8206 2488 8262 2544
rect 8206 2080 8262 2136
rect 8390 2216 8446 2272
rect 9310 8200 9366 8256
rect 9218 7928 9274 7984
rect 8852 7642 8908 7644
rect 8932 7642 8988 7644
rect 9012 7642 9068 7644
rect 9092 7642 9148 7644
rect 8852 7590 8898 7642
rect 8898 7590 8908 7642
rect 8932 7590 8962 7642
rect 8962 7590 8974 7642
rect 8974 7590 8988 7642
rect 9012 7590 9026 7642
rect 9026 7590 9038 7642
rect 9038 7590 9068 7642
rect 9092 7590 9102 7642
rect 9102 7590 9148 7642
rect 8852 7588 8908 7590
rect 8932 7588 8988 7590
rect 9012 7588 9068 7590
rect 9092 7588 9148 7590
rect 9586 11192 9642 11248
rect 9770 12144 9826 12200
rect 9678 10920 9734 10976
rect 9586 9716 9642 9752
rect 9586 9696 9588 9716
rect 9588 9696 9640 9716
rect 9640 9696 9642 9716
rect 9586 9152 9642 9208
rect 9586 8628 9642 8664
rect 9586 8608 9588 8628
rect 9588 8608 9640 8628
rect 9640 8608 9642 8628
rect 8666 6976 8722 7032
rect 9126 7112 9182 7168
rect 8852 6554 8908 6556
rect 8932 6554 8988 6556
rect 9012 6554 9068 6556
rect 9092 6554 9148 6556
rect 8852 6502 8898 6554
rect 8898 6502 8908 6554
rect 8932 6502 8962 6554
rect 8962 6502 8974 6554
rect 8974 6502 8988 6554
rect 9012 6502 9026 6554
rect 9026 6502 9038 6554
rect 9038 6502 9068 6554
rect 9092 6502 9102 6554
rect 9102 6502 9148 6554
rect 8852 6500 8908 6502
rect 8932 6500 8988 6502
rect 9012 6500 9068 6502
rect 9092 6500 9148 6502
rect 8666 6296 8722 6352
rect 8850 5888 8906 5944
rect 9402 6160 9458 6216
rect 9770 10376 9826 10432
rect 9862 7792 9918 7848
rect 9862 7384 9918 7440
rect 9770 7112 9826 7168
rect 9770 6976 9826 7032
rect 9586 6604 9588 6624
rect 9588 6604 9640 6624
rect 9640 6604 9642 6624
rect 9586 6568 9642 6604
rect 10322 15272 10378 15328
rect 12800 20698 12856 20700
rect 12880 20698 12936 20700
rect 12960 20698 13016 20700
rect 13040 20698 13096 20700
rect 12800 20646 12846 20698
rect 12846 20646 12856 20698
rect 12880 20646 12910 20698
rect 12910 20646 12922 20698
rect 12922 20646 12936 20698
rect 12960 20646 12974 20698
rect 12974 20646 12986 20698
rect 12986 20646 13016 20698
rect 13040 20646 13050 20698
rect 13050 20646 13096 20698
rect 12800 20644 12856 20646
rect 12880 20644 12936 20646
rect 12960 20644 13016 20646
rect 13040 20644 13096 20646
rect 10826 20154 10882 20156
rect 10906 20154 10962 20156
rect 10986 20154 11042 20156
rect 11066 20154 11122 20156
rect 10826 20102 10872 20154
rect 10872 20102 10882 20154
rect 10906 20102 10936 20154
rect 10936 20102 10948 20154
rect 10948 20102 10962 20154
rect 10986 20102 11000 20154
rect 11000 20102 11012 20154
rect 11012 20102 11042 20154
rect 11066 20102 11076 20154
rect 11076 20102 11122 20154
rect 10826 20100 10882 20102
rect 10906 20100 10962 20102
rect 10986 20100 11042 20102
rect 11066 20100 11122 20102
rect 10826 19066 10882 19068
rect 10906 19066 10962 19068
rect 10986 19066 11042 19068
rect 11066 19066 11122 19068
rect 10826 19014 10872 19066
rect 10872 19014 10882 19066
rect 10906 19014 10936 19066
rect 10936 19014 10948 19066
rect 10948 19014 10962 19066
rect 10986 19014 11000 19066
rect 11000 19014 11012 19066
rect 11012 19014 11042 19066
rect 11066 19014 11076 19066
rect 11076 19014 11122 19066
rect 10826 19012 10882 19014
rect 10906 19012 10962 19014
rect 10986 19012 11042 19014
rect 11066 19012 11122 19014
rect 12070 18536 12126 18592
rect 10782 18400 10838 18456
rect 10826 17978 10882 17980
rect 10906 17978 10962 17980
rect 10986 17978 11042 17980
rect 11066 17978 11122 17980
rect 10826 17926 10872 17978
rect 10872 17926 10882 17978
rect 10906 17926 10936 17978
rect 10936 17926 10948 17978
rect 10948 17926 10962 17978
rect 10986 17926 11000 17978
rect 11000 17926 11012 17978
rect 11012 17926 11042 17978
rect 11066 17926 11076 17978
rect 11076 17926 11122 17978
rect 10826 17924 10882 17926
rect 10906 17924 10962 17926
rect 10986 17924 11042 17926
rect 11066 17924 11122 17926
rect 11518 17720 11574 17776
rect 11150 17584 11206 17640
rect 10690 16904 10746 16960
rect 10826 16890 10882 16892
rect 10906 16890 10962 16892
rect 10986 16890 11042 16892
rect 11066 16890 11122 16892
rect 10826 16838 10872 16890
rect 10872 16838 10882 16890
rect 10906 16838 10936 16890
rect 10936 16838 10948 16890
rect 10948 16838 10962 16890
rect 10986 16838 11000 16890
rect 11000 16838 11012 16890
rect 11012 16838 11042 16890
rect 11066 16838 11076 16890
rect 11076 16838 11122 16890
rect 10826 16836 10882 16838
rect 10906 16836 10962 16838
rect 10986 16836 11042 16838
rect 11066 16836 11122 16838
rect 10598 16768 10654 16824
rect 10598 16496 10654 16552
rect 10506 16360 10562 16416
rect 10598 15816 10654 15872
rect 10598 15680 10654 15736
rect 10506 15020 10562 15056
rect 10506 15000 10508 15020
rect 10508 15000 10560 15020
rect 10560 15000 10562 15020
rect 10506 14592 10562 14648
rect 10826 15802 10882 15804
rect 10906 15802 10962 15804
rect 10986 15802 11042 15804
rect 11066 15802 11122 15804
rect 10826 15750 10872 15802
rect 10872 15750 10882 15802
rect 10906 15750 10936 15802
rect 10936 15750 10948 15802
rect 10948 15750 10962 15802
rect 10986 15750 11000 15802
rect 11000 15750 11012 15802
rect 11012 15750 11042 15802
rect 11066 15750 11076 15802
rect 11076 15750 11122 15802
rect 10826 15748 10882 15750
rect 10906 15748 10962 15750
rect 10986 15748 11042 15750
rect 11066 15748 11122 15750
rect 10782 15544 10838 15600
rect 10966 15580 10968 15600
rect 10968 15580 11020 15600
rect 11020 15580 11022 15600
rect 10966 15544 11022 15580
rect 11058 15136 11114 15192
rect 10826 14714 10882 14716
rect 10906 14714 10962 14716
rect 10986 14714 11042 14716
rect 11066 14714 11122 14716
rect 10826 14662 10872 14714
rect 10872 14662 10882 14714
rect 10906 14662 10936 14714
rect 10936 14662 10948 14714
rect 10948 14662 10962 14714
rect 10986 14662 11000 14714
rect 11000 14662 11012 14714
rect 11012 14662 11042 14714
rect 11066 14662 11076 14714
rect 11076 14662 11122 14714
rect 10826 14660 10882 14662
rect 10906 14660 10962 14662
rect 10986 14660 11042 14662
rect 11066 14660 11122 14662
rect 10782 14456 10838 14512
rect 10966 14456 11022 14512
rect 10230 12552 10286 12608
rect 10138 12280 10194 12336
rect 10230 12008 10286 12064
rect 10230 11872 10286 11928
rect 11702 16632 11758 16688
rect 11702 16224 11758 16280
rect 11518 15852 11520 15872
rect 11520 15852 11572 15872
rect 11572 15852 11574 15872
rect 11518 15816 11574 15852
rect 11702 15680 11758 15736
rect 11610 15000 11666 15056
rect 10826 13626 10882 13628
rect 10906 13626 10962 13628
rect 10986 13626 11042 13628
rect 11066 13626 11122 13628
rect 10826 13574 10872 13626
rect 10872 13574 10882 13626
rect 10906 13574 10936 13626
rect 10936 13574 10948 13626
rect 10948 13574 10962 13626
rect 10986 13574 11000 13626
rect 11000 13574 11012 13626
rect 11012 13574 11042 13626
rect 11066 13574 11076 13626
rect 11076 13574 11122 13626
rect 10826 13572 10882 13574
rect 10906 13572 10962 13574
rect 10986 13572 11042 13574
rect 11066 13572 11122 13574
rect 10826 12538 10882 12540
rect 10906 12538 10962 12540
rect 10986 12538 11042 12540
rect 11066 12538 11122 12540
rect 10826 12486 10872 12538
rect 10872 12486 10882 12538
rect 10906 12486 10936 12538
rect 10936 12486 10948 12538
rect 10948 12486 10962 12538
rect 10986 12486 11000 12538
rect 11000 12486 11012 12538
rect 11012 12486 11042 12538
rect 11066 12486 11076 12538
rect 11076 12486 11122 12538
rect 10826 12484 10882 12486
rect 10906 12484 10962 12486
rect 10986 12484 11042 12486
rect 11066 12484 11122 12486
rect 10598 12008 10654 12064
rect 10138 10668 10194 10704
rect 10138 10648 10140 10668
rect 10140 10648 10192 10668
rect 10192 10648 10194 10668
rect 10046 6976 10102 7032
rect 9954 6704 10010 6760
rect 9954 6432 10010 6488
rect 9218 5888 9274 5944
rect 8942 5752 8998 5808
rect 9310 5636 9366 5672
rect 9310 5616 9312 5636
rect 9312 5616 9364 5636
rect 9364 5616 9366 5636
rect 8852 5466 8908 5468
rect 8932 5466 8988 5468
rect 9012 5466 9068 5468
rect 9092 5466 9148 5468
rect 8852 5414 8898 5466
rect 8898 5414 8908 5466
rect 8932 5414 8962 5466
rect 8962 5414 8974 5466
rect 8974 5414 8988 5466
rect 9012 5414 9026 5466
rect 9026 5414 9038 5466
rect 9038 5414 9068 5466
rect 9092 5414 9102 5466
rect 9102 5414 9148 5466
rect 8852 5412 8908 5414
rect 8932 5412 8988 5414
rect 9012 5412 9068 5414
rect 9092 5412 9148 5414
rect 8758 5072 8814 5128
rect 8850 4800 8906 4856
rect 8852 4378 8908 4380
rect 8932 4378 8988 4380
rect 9012 4378 9068 4380
rect 9092 4378 9148 4380
rect 8852 4326 8898 4378
rect 8898 4326 8908 4378
rect 8932 4326 8962 4378
rect 8962 4326 8974 4378
rect 8974 4326 8988 4378
rect 9012 4326 9026 4378
rect 9026 4326 9038 4378
rect 9038 4326 9068 4378
rect 9092 4326 9102 4378
rect 9102 4326 9148 4378
rect 8852 4324 8908 4326
rect 8932 4324 8988 4326
rect 9012 4324 9068 4326
rect 9092 4324 9148 4326
rect 9310 4256 9366 4312
rect 9494 5208 9550 5264
rect 9770 5888 9826 5944
rect 9586 5072 9642 5128
rect 11058 12280 11114 12336
rect 10966 11872 11022 11928
rect 10874 11600 10930 11656
rect 11058 11600 11114 11656
rect 10826 11450 10882 11452
rect 10906 11450 10962 11452
rect 10986 11450 11042 11452
rect 11066 11450 11122 11452
rect 10826 11398 10872 11450
rect 10872 11398 10882 11450
rect 10906 11398 10936 11450
rect 10936 11398 10948 11450
rect 10948 11398 10962 11450
rect 10986 11398 11000 11450
rect 11000 11398 11012 11450
rect 11012 11398 11042 11450
rect 11066 11398 11076 11450
rect 11076 11398 11122 11450
rect 10826 11396 10882 11398
rect 10906 11396 10962 11398
rect 10986 11396 11042 11398
rect 11066 11396 11122 11398
rect 10598 11056 10654 11112
rect 10598 10784 10654 10840
rect 10966 10920 11022 10976
rect 11334 13524 11390 13560
rect 11334 13504 11336 13524
rect 11336 13504 11388 13524
rect 11388 13504 11390 13524
rect 11426 13096 11482 13152
rect 11334 12960 11390 13016
rect 11886 14456 11942 14512
rect 11610 14048 11666 14104
rect 11794 14048 11850 14104
rect 11518 12960 11574 13016
rect 11518 12552 11574 12608
rect 10826 10362 10882 10364
rect 10906 10362 10962 10364
rect 10986 10362 11042 10364
rect 11066 10362 11122 10364
rect 10826 10310 10872 10362
rect 10872 10310 10882 10362
rect 10906 10310 10936 10362
rect 10936 10310 10948 10362
rect 10948 10310 10962 10362
rect 10986 10310 11000 10362
rect 11000 10310 11012 10362
rect 11012 10310 11042 10362
rect 11066 10310 11076 10362
rect 11076 10310 11122 10362
rect 10826 10308 10882 10310
rect 10906 10308 10962 10310
rect 10986 10308 11042 10310
rect 11066 10308 11122 10310
rect 10690 9424 10746 9480
rect 10826 9274 10882 9276
rect 10906 9274 10962 9276
rect 10986 9274 11042 9276
rect 11066 9274 11122 9276
rect 10826 9222 10872 9274
rect 10872 9222 10882 9274
rect 10906 9222 10936 9274
rect 10936 9222 10948 9274
rect 10948 9222 10962 9274
rect 10986 9222 11000 9274
rect 11000 9222 11012 9274
rect 11012 9222 11042 9274
rect 11066 9222 11076 9274
rect 11076 9222 11122 9274
rect 10826 9220 10882 9222
rect 10906 9220 10962 9222
rect 10986 9220 11042 9222
rect 11066 9220 11122 9222
rect 11794 12416 11850 12472
rect 11702 11872 11758 11928
rect 11426 11192 11482 11248
rect 11334 10376 11390 10432
rect 11242 10240 11298 10296
rect 10874 8608 10930 8664
rect 10826 8186 10882 8188
rect 10906 8186 10962 8188
rect 10986 8186 11042 8188
rect 11066 8186 11122 8188
rect 10826 8134 10872 8186
rect 10872 8134 10882 8186
rect 10906 8134 10936 8186
rect 10936 8134 10948 8186
rect 10948 8134 10962 8186
rect 10986 8134 11000 8186
rect 11000 8134 11012 8186
rect 11012 8134 11042 8186
rect 11066 8134 11076 8186
rect 11076 8134 11122 8186
rect 10826 8132 10882 8134
rect 10906 8132 10962 8134
rect 10986 8132 11042 8134
rect 11066 8132 11122 8134
rect 10782 7928 10838 7984
rect 10966 7792 11022 7848
rect 10966 7384 11022 7440
rect 10414 6160 10470 6216
rect 10322 6060 10324 6080
rect 10324 6060 10376 6080
rect 10376 6060 10378 6080
rect 10322 6024 10378 6060
rect 10230 5788 10232 5808
rect 10232 5788 10284 5808
rect 10284 5788 10286 5808
rect 10230 5752 10286 5788
rect 9770 5208 9826 5264
rect 9678 4800 9734 4856
rect 9678 4664 9734 4720
rect 9126 3712 9182 3768
rect 9310 3304 9366 3360
rect 8852 3290 8908 3292
rect 8932 3290 8988 3292
rect 9012 3290 9068 3292
rect 9092 3290 9148 3292
rect 8852 3238 8898 3290
rect 8898 3238 8908 3290
rect 8932 3238 8962 3290
rect 8962 3238 8974 3290
rect 8974 3238 8988 3290
rect 9012 3238 9026 3290
rect 9026 3238 9038 3290
rect 9038 3238 9068 3290
rect 9092 3238 9102 3290
rect 9102 3238 9148 3290
rect 8852 3236 8908 3238
rect 8932 3236 8988 3238
rect 9012 3236 9068 3238
rect 9092 3236 9148 3238
rect 8758 2352 8814 2408
rect 9310 3168 9366 3224
rect 9402 3032 9458 3088
rect 8852 2202 8908 2204
rect 8932 2202 8988 2204
rect 9012 2202 9068 2204
rect 9092 2202 9148 2204
rect 8852 2150 8898 2202
rect 8898 2150 8908 2202
rect 8932 2150 8962 2202
rect 8962 2150 8974 2202
rect 8974 2150 8988 2202
rect 9012 2150 9026 2202
rect 9026 2150 9038 2202
rect 9038 2150 9068 2202
rect 9092 2150 9102 2202
rect 9102 2150 9148 2202
rect 8852 2148 8908 2150
rect 8932 2148 8988 2150
rect 9012 2148 9068 2150
rect 9092 2148 9148 2150
rect 8758 1264 8814 1320
rect 9310 2216 9366 2272
rect 9218 1400 9274 1456
rect 8574 1128 8630 1184
rect 8852 1114 8908 1116
rect 8932 1114 8988 1116
rect 9012 1114 9068 1116
rect 9092 1114 9148 1116
rect 8852 1062 8898 1114
rect 8898 1062 8908 1114
rect 8932 1062 8962 1114
rect 8962 1062 8974 1114
rect 8974 1062 8988 1114
rect 9012 1062 9026 1114
rect 9026 1062 9038 1114
rect 9038 1062 9068 1114
rect 9092 1062 9102 1114
rect 9102 1062 9148 1114
rect 8852 1060 8908 1062
rect 8932 1060 8988 1062
rect 9012 1060 9068 1062
rect 9092 1060 9148 1062
rect 7930 720 7986 776
rect 8206 720 8262 776
rect 9494 992 9550 1048
rect 10506 5888 10562 5944
rect 10506 5616 10562 5672
rect 10826 7098 10882 7100
rect 10906 7098 10962 7100
rect 10986 7098 11042 7100
rect 11066 7098 11122 7100
rect 10826 7046 10872 7098
rect 10872 7046 10882 7098
rect 10906 7046 10936 7098
rect 10936 7046 10948 7098
rect 10948 7046 10962 7098
rect 10986 7046 11000 7098
rect 11000 7046 11012 7098
rect 11012 7046 11042 7098
rect 11066 7046 11076 7098
rect 11076 7046 11122 7098
rect 10826 7044 10882 7046
rect 10906 7044 10962 7046
rect 10986 7044 11042 7046
rect 11066 7044 11122 7046
rect 11058 6840 11114 6896
rect 10598 5480 10654 5536
rect 10230 4664 10286 4720
rect 10874 6568 10930 6624
rect 11058 6568 11114 6624
rect 11334 9152 11390 9208
rect 11702 11464 11758 11520
rect 11242 8200 11298 8256
rect 11426 7792 11482 7848
rect 11242 6976 11298 7032
rect 11058 6296 11114 6352
rect 10826 6010 10882 6012
rect 10906 6010 10962 6012
rect 10986 6010 11042 6012
rect 11066 6010 11122 6012
rect 10826 5958 10872 6010
rect 10872 5958 10882 6010
rect 10906 5958 10936 6010
rect 10936 5958 10948 6010
rect 10948 5958 10962 6010
rect 10986 5958 11000 6010
rect 11000 5958 11012 6010
rect 11012 5958 11042 6010
rect 11066 5958 11076 6010
rect 11076 5958 11122 6010
rect 10826 5956 10882 5958
rect 10906 5956 10962 5958
rect 10986 5956 11042 5958
rect 11066 5956 11122 5958
rect 11058 5752 11114 5808
rect 10782 5616 10838 5672
rect 10826 4922 10882 4924
rect 10906 4922 10962 4924
rect 10986 4922 11042 4924
rect 11066 4922 11122 4924
rect 10826 4870 10872 4922
rect 10872 4870 10882 4922
rect 10906 4870 10936 4922
rect 10936 4870 10948 4922
rect 10948 4870 10962 4922
rect 10986 4870 11000 4922
rect 11000 4870 11012 4922
rect 11012 4870 11042 4922
rect 11066 4870 11076 4922
rect 11076 4870 11122 4922
rect 10826 4868 10882 4870
rect 10906 4868 10962 4870
rect 10986 4868 11042 4870
rect 11066 4868 11122 4870
rect 10598 4800 10654 4856
rect 10230 3168 10286 3224
rect 10230 2760 10286 2816
rect 9862 2080 9918 2136
rect 10138 1808 10194 1864
rect 10230 1536 10286 1592
rect 9954 1264 10010 1320
rect 9678 448 9734 504
rect 10690 4256 10746 4312
rect 10506 3848 10562 3904
rect 11242 4256 11298 4312
rect 10826 3834 10882 3836
rect 10906 3834 10962 3836
rect 10986 3834 11042 3836
rect 11066 3834 11122 3836
rect 10826 3782 10872 3834
rect 10872 3782 10882 3834
rect 10906 3782 10936 3834
rect 10936 3782 10948 3834
rect 10948 3782 10962 3834
rect 10986 3782 11000 3834
rect 11000 3782 11012 3834
rect 11012 3782 11042 3834
rect 11066 3782 11076 3834
rect 11076 3782 11122 3834
rect 10826 3780 10882 3782
rect 10906 3780 10962 3782
rect 10986 3780 11042 3782
rect 11066 3780 11122 3782
rect 10966 3032 11022 3088
rect 11242 3848 11298 3904
rect 10826 2746 10882 2748
rect 10906 2746 10962 2748
rect 10986 2746 11042 2748
rect 11066 2746 11122 2748
rect 10826 2694 10872 2746
rect 10872 2694 10882 2746
rect 10906 2694 10936 2746
rect 10936 2694 10948 2746
rect 10948 2694 10962 2746
rect 10986 2694 11000 2746
rect 11000 2694 11012 2746
rect 11012 2694 11042 2746
rect 11066 2694 11076 2746
rect 11076 2694 11122 2746
rect 10826 2692 10882 2694
rect 10906 2692 10962 2694
rect 10986 2692 11042 2694
rect 11066 2692 11122 2694
rect 10874 2488 10930 2544
rect 10782 2080 10838 2136
rect 10874 1808 10930 1864
rect 10826 1658 10882 1660
rect 10906 1658 10962 1660
rect 10986 1658 11042 1660
rect 11066 1658 11122 1660
rect 10826 1606 10872 1658
rect 10872 1606 10882 1658
rect 10906 1606 10936 1658
rect 10936 1606 10948 1658
rect 10948 1606 10962 1658
rect 10986 1606 11000 1658
rect 11000 1606 11012 1658
rect 11012 1606 11042 1658
rect 11066 1606 11076 1658
rect 11076 1606 11122 1658
rect 10826 1604 10882 1606
rect 10906 1604 10962 1606
rect 10986 1604 11042 1606
rect 11066 1604 11122 1606
rect 11610 7268 11666 7304
rect 11610 7248 11612 7268
rect 11612 7248 11664 7268
rect 11664 7248 11666 7268
rect 11610 6296 11666 6352
rect 11610 5888 11666 5944
rect 11610 4936 11666 4992
rect 12346 17176 12402 17232
rect 12162 15272 12218 15328
rect 12070 15136 12126 15192
rect 12070 14864 12126 14920
rect 12800 19610 12856 19612
rect 12880 19610 12936 19612
rect 12960 19610 13016 19612
rect 13040 19610 13096 19612
rect 12800 19558 12846 19610
rect 12846 19558 12856 19610
rect 12880 19558 12910 19610
rect 12910 19558 12922 19610
rect 12922 19558 12936 19610
rect 12960 19558 12974 19610
rect 12974 19558 12986 19610
rect 12986 19558 13016 19610
rect 13040 19558 13050 19610
rect 13050 19558 13096 19610
rect 12800 19556 12856 19558
rect 12880 19556 12936 19558
rect 12960 19556 13016 19558
rect 13040 19556 13096 19558
rect 12800 18522 12856 18524
rect 12880 18522 12936 18524
rect 12960 18522 13016 18524
rect 13040 18522 13096 18524
rect 12800 18470 12846 18522
rect 12846 18470 12856 18522
rect 12880 18470 12910 18522
rect 12910 18470 12922 18522
rect 12922 18470 12936 18522
rect 12960 18470 12974 18522
rect 12974 18470 12986 18522
rect 12986 18470 13016 18522
rect 13040 18470 13050 18522
rect 13050 18470 13096 18522
rect 12800 18468 12856 18470
rect 12880 18468 12936 18470
rect 12960 18468 13016 18470
rect 13040 18468 13096 18470
rect 12800 17434 12856 17436
rect 12880 17434 12936 17436
rect 12960 17434 13016 17436
rect 13040 17434 13096 17436
rect 12800 17382 12846 17434
rect 12846 17382 12856 17434
rect 12880 17382 12910 17434
rect 12910 17382 12922 17434
rect 12922 17382 12936 17434
rect 12960 17382 12974 17434
rect 12974 17382 12986 17434
rect 12986 17382 13016 17434
rect 13040 17382 13050 17434
rect 13050 17382 13096 17434
rect 12800 17380 12856 17382
rect 12880 17380 12936 17382
rect 12960 17380 13016 17382
rect 13040 17380 13096 17382
rect 12800 16346 12856 16348
rect 12880 16346 12936 16348
rect 12960 16346 13016 16348
rect 13040 16346 13096 16348
rect 12800 16294 12846 16346
rect 12846 16294 12856 16346
rect 12880 16294 12910 16346
rect 12910 16294 12922 16346
rect 12922 16294 12936 16346
rect 12960 16294 12974 16346
rect 12974 16294 12986 16346
rect 12986 16294 13016 16346
rect 13040 16294 13050 16346
rect 13050 16294 13096 16346
rect 12800 16292 12856 16294
rect 12880 16292 12936 16294
rect 12960 16292 13016 16294
rect 13040 16292 13096 16294
rect 13082 16088 13138 16144
rect 12162 14184 12218 14240
rect 12070 14048 12126 14104
rect 12070 13640 12126 13696
rect 12162 13232 12218 13288
rect 13174 15816 13230 15872
rect 12898 15564 12954 15600
rect 12898 15544 12900 15564
rect 12900 15544 12952 15564
rect 12952 15544 12954 15564
rect 12714 15408 12770 15464
rect 12990 15444 12992 15464
rect 12992 15444 13044 15464
rect 13044 15444 13046 15464
rect 12990 15408 13046 15444
rect 12070 11756 12126 11792
rect 12070 11736 12072 11756
rect 12072 11736 12124 11756
rect 12124 11736 12126 11756
rect 12254 12416 12310 12472
rect 12254 12008 12310 12064
rect 12622 14864 12678 14920
rect 12530 13268 12532 13288
rect 12532 13268 12584 13288
rect 12584 13268 12586 13288
rect 12530 13232 12586 13268
rect 12438 13096 12494 13152
rect 12438 12960 12494 13016
rect 12438 12688 12494 12744
rect 12346 11872 12402 11928
rect 12254 11328 12310 11384
rect 12800 15258 12856 15260
rect 12880 15258 12936 15260
rect 12960 15258 13016 15260
rect 13040 15258 13096 15260
rect 12800 15206 12846 15258
rect 12846 15206 12856 15258
rect 12880 15206 12910 15258
rect 12910 15206 12922 15258
rect 12922 15206 12936 15258
rect 12960 15206 12974 15258
rect 12974 15206 12986 15258
rect 12986 15206 13016 15258
rect 13040 15206 13050 15258
rect 13050 15206 13096 15258
rect 12800 15204 12856 15206
rect 12880 15204 12936 15206
rect 12960 15204 13016 15206
rect 13040 15204 13096 15206
rect 12714 14592 12770 14648
rect 12800 14170 12856 14172
rect 12880 14170 12936 14172
rect 12960 14170 13016 14172
rect 13040 14170 13096 14172
rect 12800 14118 12846 14170
rect 12846 14118 12856 14170
rect 12880 14118 12910 14170
rect 12910 14118 12922 14170
rect 12922 14118 12936 14170
rect 12960 14118 12974 14170
rect 12974 14118 12986 14170
rect 12986 14118 13016 14170
rect 13040 14118 13050 14170
rect 13050 14118 13096 14170
rect 12800 14116 12856 14118
rect 12880 14116 12936 14118
rect 12960 14116 13016 14118
rect 13040 14116 13096 14118
rect 12714 13776 12770 13832
rect 12990 13504 13046 13560
rect 12800 13082 12856 13084
rect 12880 13082 12936 13084
rect 12960 13082 13016 13084
rect 13040 13082 13096 13084
rect 12800 13030 12846 13082
rect 12846 13030 12856 13082
rect 12880 13030 12910 13082
rect 12910 13030 12922 13082
rect 12922 13030 12936 13082
rect 12960 13030 12974 13082
rect 12974 13030 12986 13082
rect 12986 13030 13016 13082
rect 13040 13030 13050 13082
rect 13050 13030 13096 13082
rect 12800 13028 12856 13030
rect 12880 13028 12936 13030
rect 12960 13028 13016 13030
rect 13040 13028 13096 13030
rect 12898 12688 12954 12744
rect 13174 12436 13230 12472
rect 13174 12416 13176 12436
rect 13176 12416 13228 12436
rect 13228 12416 13230 12436
rect 13542 14728 13598 14784
rect 13542 14476 13598 14512
rect 13542 14456 13544 14476
rect 13544 14456 13596 14476
rect 13596 14456 13598 14476
rect 13726 15544 13782 15600
rect 13450 14184 13506 14240
rect 13450 13776 13506 13832
rect 13542 13504 13598 13560
rect 13450 12960 13506 13016
rect 13726 13504 13782 13560
rect 12800 11994 12856 11996
rect 12880 11994 12936 11996
rect 12960 11994 13016 11996
rect 13040 11994 13096 11996
rect 12800 11942 12846 11994
rect 12846 11942 12856 11994
rect 12880 11942 12910 11994
rect 12910 11942 12922 11994
rect 12922 11942 12936 11994
rect 12960 11942 12974 11994
rect 12974 11942 12986 11994
rect 12986 11942 13016 11994
rect 13040 11942 13050 11994
rect 13050 11942 13096 11994
rect 12800 11940 12856 11942
rect 12880 11940 12936 11942
rect 12960 11940 13016 11942
rect 13040 11940 13096 11942
rect 12530 11328 12586 11384
rect 12162 11092 12164 11112
rect 12164 11092 12216 11112
rect 12216 11092 12218 11112
rect 12162 11056 12218 11092
rect 11794 9560 11850 9616
rect 11978 9696 12034 9752
rect 11978 9596 11980 9616
rect 11980 9596 12032 9616
rect 12032 9596 12034 9616
rect 11978 9560 12034 9596
rect 11886 7792 11942 7848
rect 12254 10784 12310 10840
rect 11978 6432 12034 6488
rect 11886 5772 11942 5808
rect 11886 5752 11888 5772
rect 11888 5752 11940 5772
rect 11940 5752 11942 5772
rect 12530 9832 12586 9888
rect 12346 9288 12402 9344
rect 12530 8880 12586 8936
rect 12530 8608 12586 8664
rect 12438 7792 12494 7848
rect 12438 7656 12494 7712
rect 12438 7112 12494 7168
rect 11886 5480 11942 5536
rect 11886 5344 11942 5400
rect 12162 5344 12218 5400
rect 12162 5072 12218 5128
rect 13450 12316 13452 12336
rect 13452 12316 13504 12336
rect 13504 12316 13506 12336
rect 14002 14068 14058 14104
rect 14002 14048 14004 14068
rect 14004 14048 14056 14068
rect 14056 14048 14058 14068
rect 14002 13912 14058 13968
rect 13910 13776 13966 13832
rect 13818 12824 13874 12880
rect 13450 12280 13506 12316
rect 13450 11872 13506 11928
rect 13726 12008 13782 12064
rect 14002 13640 14058 13696
rect 14186 13640 14242 13696
rect 14186 12960 14242 13016
rect 14186 12688 14242 12744
rect 14002 12552 14058 12608
rect 14094 12300 14150 12336
rect 14094 12280 14096 12300
rect 14096 12280 14148 12300
rect 14148 12280 14150 12300
rect 13726 11464 13782 11520
rect 12800 10906 12856 10908
rect 12880 10906 12936 10908
rect 12960 10906 13016 10908
rect 13040 10906 13096 10908
rect 12800 10854 12846 10906
rect 12846 10854 12856 10906
rect 12880 10854 12910 10906
rect 12910 10854 12922 10906
rect 12922 10854 12936 10906
rect 12960 10854 12974 10906
rect 12974 10854 12986 10906
rect 12986 10854 13016 10906
rect 13040 10854 13050 10906
rect 13050 10854 13096 10906
rect 12800 10852 12856 10854
rect 12880 10852 12936 10854
rect 12960 10852 13016 10854
rect 13040 10852 13096 10854
rect 13266 10920 13322 10976
rect 12806 10512 12862 10568
rect 13174 10512 13230 10568
rect 13358 10376 13414 10432
rect 12990 10004 12992 10024
rect 12992 10004 13044 10024
rect 13044 10004 13046 10024
rect 12990 9968 13046 10004
rect 12800 9818 12856 9820
rect 12880 9818 12936 9820
rect 12960 9818 13016 9820
rect 13040 9818 13096 9820
rect 12800 9766 12846 9818
rect 12846 9766 12856 9818
rect 12880 9766 12910 9818
rect 12910 9766 12922 9818
rect 12922 9766 12936 9818
rect 12960 9766 12974 9818
rect 12974 9766 12986 9818
rect 12986 9766 13016 9818
rect 13040 9766 13050 9818
rect 13050 9766 13096 9818
rect 12800 9764 12856 9766
rect 12880 9764 12936 9766
rect 12960 9764 13016 9766
rect 13040 9764 13096 9766
rect 12990 8916 12992 8936
rect 12992 8916 13044 8936
rect 13044 8916 13046 8936
rect 12990 8880 13046 8916
rect 13450 10240 13506 10296
rect 13450 9832 13506 9888
rect 13266 9016 13322 9072
rect 12800 8730 12856 8732
rect 12880 8730 12936 8732
rect 12960 8730 13016 8732
rect 13040 8730 13096 8732
rect 12800 8678 12846 8730
rect 12846 8678 12856 8730
rect 12880 8678 12910 8730
rect 12910 8678 12922 8730
rect 12922 8678 12936 8730
rect 12960 8678 12974 8730
rect 12974 8678 12986 8730
rect 12986 8678 13016 8730
rect 13040 8678 13050 8730
rect 13050 8678 13096 8730
rect 12800 8676 12856 8678
rect 12880 8676 12936 8678
rect 12960 8676 13016 8678
rect 13040 8676 13096 8678
rect 12714 7928 12770 7984
rect 12898 7928 12954 7984
rect 12800 7642 12856 7644
rect 12880 7642 12936 7644
rect 12960 7642 13016 7644
rect 13040 7642 13096 7644
rect 12800 7590 12846 7642
rect 12846 7590 12856 7642
rect 12880 7590 12910 7642
rect 12910 7590 12922 7642
rect 12922 7590 12936 7642
rect 12960 7590 12974 7642
rect 12974 7590 12986 7642
rect 12986 7590 13016 7642
rect 13040 7590 13050 7642
rect 13050 7590 13096 7642
rect 12800 7588 12856 7590
rect 12880 7588 12936 7590
rect 12960 7588 13016 7590
rect 13040 7588 13096 7590
rect 13634 9424 13690 9480
rect 14002 10920 14058 10976
rect 13910 10376 13966 10432
rect 13726 8608 13782 8664
rect 13726 8508 13728 8528
rect 13728 8508 13780 8528
rect 13780 8508 13782 8528
rect 13726 8472 13782 8508
rect 12622 6568 12678 6624
rect 12800 6554 12856 6556
rect 12880 6554 12936 6556
rect 12960 6554 13016 6556
rect 13040 6554 13096 6556
rect 12800 6502 12846 6554
rect 12846 6502 12856 6554
rect 12880 6502 12910 6554
rect 12910 6502 12922 6554
rect 12922 6502 12936 6554
rect 12960 6502 12974 6554
rect 12974 6502 12986 6554
rect 12986 6502 13016 6554
rect 13040 6502 13050 6554
rect 13050 6502 13096 6554
rect 12800 6500 12856 6502
rect 12880 6500 12936 6502
rect 12960 6500 13016 6502
rect 13040 6500 13096 6502
rect 12806 6296 12862 6352
rect 12530 5344 12586 5400
rect 12346 5092 12402 5128
rect 12346 5072 12348 5092
rect 12348 5072 12400 5092
rect 12400 5072 12402 5092
rect 12622 4936 12678 4992
rect 11978 4528 12034 4584
rect 11886 4256 11942 4312
rect 11702 3612 11704 3632
rect 11704 3612 11756 3632
rect 11756 3612 11758 3632
rect 11702 3576 11758 3612
rect 12070 4392 12126 4448
rect 11886 3304 11942 3360
rect 12346 4140 12402 4176
rect 12346 4120 12348 4140
rect 12348 4120 12400 4140
rect 12400 4120 12402 4140
rect 11702 3032 11758 3088
rect 11334 1672 11390 1728
rect 12070 2624 12126 2680
rect 12162 2352 12218 2408
rect 12622 4256 12678 4312
rect 12622 3848 12678 3904
rect 13450 6840 13506 6896
rect 13266 6568 13322 6624
rect 13174 5752 13230 5808
rect 12800 5466 12856 5468
rect 12880 5466 12936 5468
rect 12960 5466 13016 5468
rect 13040 5466 13096 5468
rect 12800 5414 12846 5466
rect 12846 5414 12856 5466
rect 12880 5414 12910 5466
rect 12910 5414 12922 5466
rect 12922 5414 12936 5466
rect 12960 5414 12974 5466
rect 12974 5414 12986 5466
rect 12986 5414 13016 5466
rect 13040 5414 13050 5466
rect 13050 5414 13096 5466
rect 12800 5412 12856 5414
rect 12880 5412 12936 5414
rect 12960 5412 13016 5414
rect 13040 5412 13096 5414
rect 12806 4800 12862 4856
rect 13542 6432 13598 6488
rect 13358 5752 13414 5808
rect 12800 4378 12856 4380
rect 12880 4378 12936 4380
rect 12960 4378 13016 4380
rect 13040 4378 13096 4380
rect 12800 4326 12846 4378
rect 12846 4326 12856 4378
rect 12880 4326 12910 4378
rect 12910 4326 12922 4378
rect 12922 4326 12936 4378
rect 12960 4326 12974 4378
rect 12974 4326 12986 4378
rect 12986 4326 13016 4378
rect 13040 4326 13050 4378
rect 13050 4326 13096 4378
rect 12800 4324 12856 4326
rect 12880 4324 12936 4326
rect 12960 4324 13016 4326
rect 13040 4324 13096 4326
rect 13542 4528 13598 4584
rect 14774 21242 14830 21244
rect 14854 21242 14910 21244
rect 14934 21242 14990 21244
rect 15014 21242 15070 21244
rect 14774 21190 14820 21242
rect 14820 21190 14830 21242
rect 14854 21190 14884 21242
rect 14884 21190 14896 21242
rect 14896 21190 14910 21242
rect 14934 21190 14948 21242
rect 14948 21190 14960 21242
rect 14960 21190 14990 21242
rect 15014 21190 15024 21242
rect 15024 21190 15070 21242
rect 14774 21188 14830 21190
rect 14854 21188 14910 21190
rect 14934 21188 14990 21190
rect 15014 21188 15070 21190
rect 14774 20154 14830 20156
rect 14854 20154 14910 20156
rect 14934 20154 14990 20156
rect 15014 20154 15070 20156
rect 14774 20102 14820 20154
rect 14820 20102 14830 20154
rect 14854 20102 14884 20154
rect 14884 20102 14896 20154
rect 14896 20102 14910 20154
rect 14934 20102 14948 20154
rect 14948 20102 14960 20154
rect 14960 20102 14990 20154
rect 15014 20102 15024 20154
rect 15024 20102 15070 20154
rect 14774 20100 14830 20102
rect 14854 20100 14910 20102
rect 14934 20100 14990 20102
rect 15014 20100 15070 20102
rect 14774 19066 14830 19068
rect 14854 19066 14910 19068
rect 14934 19066 14990 19068
rect 15014 19066 15070 19068
rect 14774 19014 14820 19066
rect 14820 19014 14830 19066
rect 14854 19014 14884 19066
rect 14884 19014 14896 19066
rect 14896 19014 14910 19066
rect 14934 19014 14948 19066
rect 14948 19014 14960 19066
rect 14960 19014 14990 19066
rect 15014 19014 15024 19066
rect 15024 19014 15070 19066
rect 14774 19012 14830 19014
rect 14854 19012 14910 19014
rect 14934 19012 14990 19014
rect 15014 19012 15070 19014
rect 15198 18672 15254 18728
rect 14774 17978 14830 17980
rect 14854 17978 14910 17980
rect 14934 17978 14990 17980
rect 15014 17978 15070 17980
rect 14774 17926 14820 17978
rect 14820 17926 14830 17978
rect 14854 17926 14884 17978
rect 14884 17926 14896 17978
rect 14896 17926 14910 17978
rect 14934 17926 14948 17978
rect 14948 17926 14960 17978
rect 14960 17926 14990 17978
rect 15014 17926 15024 17978
rect 15024 17926 15070 17978
rect 14774 17924 14830 17926
rect 14854 17924 14910 17926
rect 14934 17924 14990 17926
rect 15014 17924 15070 17926
rect 14774 16890 14830 16892
rect 14854 16890 14910 16892
rect 14934 16890 14990 16892
rect 15014 16890 15070 16892
rect 14774 16838 14820 16890
rect 14820 16838 14830 16890
rect 14854 16838 14884 16890
rect 14884 16838 14896 16890
rect 14896 16838 14910 16890
rect 14934 16838 14948 16890
rect 14948 16838 14960 16890
rect 14960 16838 14990 16890
rect 15014 16838 15024 16890
rect 15024 16838 15070 16890
rect 14774 16836 14830 16838
rect 14854 16836 14910 16838
rect 14934 16836 14990 16838
rect 15014 16836 15070 16838
rect 14774 15802 14830 15804
rect 14854 15802 14910 15804
rect 14934 15802 14990 15804
rect 15014 15802 15070 15804
rect 14774 15750 14820 15802
rect 14820 15750 14830 15802
rect 14854 15750 14884 15802
rect 14884 15750 14896 15802
rect 14896 15750 14910 15802
rect 14934 15750 14948 15802
rect 14948 15750 14960 15802
rect 14960 15750 14990 15802
rect 15014 15750 15024 15802
rect 15024 15750 15070 15802
rect 14774 15748 14830 15750
rect 14854 15748 14910 15750
rect 14934 15748 14990 15750
rect 15014 15748 15070 15750
rect 14774 14714 14830 14716
rect 14854 14714 14910 14716
rect 14934 14714 14990 14716
rect 15014 14714 15070 14716
rect 14774 14662 14820 14714
rect 14820 14662 14830 14714
rect 14854 14662 14884 14714
rect 14884 14662 14896 14714
rect 14896 14662 14910 14714
rect 14934 14662 14948 14714
rect 14948 14662 14960 14714
rect 14960 14662 14990 14714
rect 15014 14662 15024 14714
rect 15024 14662 15070 14714
rect 14774 14660 14830 14662
rect 14854 14660 14910 14662
rect 14934 14660 14990 14662
rect 15014 14660 15070 14662
rect 14922 14356 14924 14376
rect 14924 14356 14976 14376
rect 14976 14356 14978 14376
rect 14922 14320 14978 14356
rect 14554 13776 14610 13832
rect 14462 13640 14518 13696
rect 14370 12960 14426 13016
rect 14370 12824 14426 12880
rect 14370 12144 14426 12200
rect 14278 10376 14334 10432
rect 14186 10104 14242 10160
rect 14094 9832 14150 9888
rect 14278 9868 14280 9888
rect 14280 9868 14332 9888
rect 14332 9868 14334 9888
rect 14278 9832 14334 9868
rect 14186 9152 14242 9208
rect 14002 9016 14058 9072
rect 13910 8064 13966 8120
rect 13818 7792 13874 7848
rect 13910 7540 13966 7576
rect 13910 7520 13912 7540
rect 13912 7520 13964 7540
rect 13964 7520 13966 7540
rect 13910 7248 13966 7304
rect 13174 3848 13230 3904
rect 12806 3712 12862 3768
rect 12622 3168 12678 3224
rect 12806 3440 12862 3496
rect 12800 3290 12856 3292
rect 12880 3290 12936 3292
rect 12960 3290 13016 3292
rect 13040 3290 13096 3292
rect 12800 3238 12846 3290
rect 12846 3238 12856 3290
rect 12880 3238 12910 3290
rect 12910 3238 12922 3290
rect 12922 3238 12936 3290
rect 12960 3238 12974 3290
rect 12974 3238 12986 3290
rect 12986 3238 13016 3290
rect 13040 3238 13050 3290
rect 13050 3238 13096 3290
rect 12800 3236 12856 3238
rect 12880 3236 12936 3238
rect 12960 3236 13016 3238
rect 13040 3236 13096 3238
rect 12346 2624 12402 2680
rect 11794 1844 11796 1864
rect 11796 1844 11848 1864
rect 11848 1844 11850 1864
rect 11794 1808 11850 1844
rect 11702 1556 11758 1592
rect 11702 1536 11704 1556
rect 11704 1536 11756 1556
rect 11756 1536 11758 1556
rect 11886 584 11942 640
rect 12438 2080 12494 2136
rect 13174 2216 13230 2272
rect 12800 2202 12856 2204
rect 12880 2202 12936 2204
rect 12960 2202 13016 2204
rect 13040 2202 13096 2204
rect 12800 2150 12846 2202
rect 12846 2150 12856 2202
rect 12880 2150 12910 2202
rect 12910 2150 12922 2202
rect 12922 2150 12936 2202
rect 12960 2150 12974 2202
rect 12974 2150 12986 2202
rect 12986 2150 13016 2202
rect 13040 2150 13050 2202
rect 13050 2150 13096 2202
rect 12800 2148 12856 2150
rect 12880 2148 12936 2150
rect 12960 2148 13016 2150
rect 13040 2148 13096 2150
rect 12990 1808 13046 1864
rect 13266 1672 13322 1728
rect 12800 1114 12856 1116
rect 12880 1114 12936 1116
rect 12960 1114 13016 1116
rect 13040 1114 13096 1116
rect 12800 1062 12846 1114
rect 12846 1062 12856 1114
rect 12880 1062 12910 1114
rect 12910 1062 12922 1114
rect 12922 1062 12936 1114
rect 12960 1062 12974 1114
rect 12974 1062 12986 1114
rect 12986 1062 13016 1114
rect 13040 1062 13050 1114
rect 13050 1062 13096 1114
rect 12800 1060 12856 1062
rect 12880 1060 12936 1062
rect 12960 1060 13016 1062
rect 13040 1060 13096 1062
rect 12530 992 12586 1048
rect 13726 3984 13782 4040
rect 13726 3848 13782 3904
rect 13542 2760 13598 2816
rect 13726 3304 13782 3360
rect 14094 8064 14150 8120
rect 14186 6024 14242 6080
rect 13726 3052 13782 3088
rect 13726 3032 13728 3052
rect 13728 3032 13780 3052
rect 13780 3032 13782 3052
rect 13542 1264 13598 1320
rect 13266 448 13322 504
rect 14094 4256 14150 4312
rect 14094 3848 14150 3904
rect 14094 3068 14096 3088
rect 14096 3068 14148 3088
rect 14148 3068 14150 3088
rect 14094 3032 14150 3068
rect 14002 2624 14058 2680
rect 14278 4820 14334 4856
rect 14278 4800 14280 4820
rect 14280 4800 14332 4820
rect 14332 4800 14334 4820
rect 15106 13776 15162 13832
rect 14774 13626 14830 13628
rect 14854 13626 14910 13628
rect 14934 13626 14990 13628
rect 15014 13626 15070 13628
rect 14774 13574 14820 13626
rect 14820 13574 14830 13626
rect 14854 13574 14884 13626
rect 14884 13574 14896 13626
rect 14896 13574 14910 13626
rect 14934 13574 14948 13626
rect 14948 13574 14960 13626
rect 14960 13574 14990 13626
rect 15014 13574 15024 13626
rect 15024 13574 15070 13626
rect 14774 13572 14830 13574
rect 14854 13572 14910 13574
rect 14934 13572 14990 13574
rect 15014 13572 15070 13574
rect 14830 12688 14886 12744
rect 14774 12538 14830 12540
rect 14854 12538 14910 12540
rect 14934 12538 14990 12540
rect 15014 12538 15070 12540
rect 14774 12486 14820 12538
rect 14820 12486 14830 12538
rect 14854 12486 14884 12538
rect 14884 12486 14896 12538
rect 14896 12486 14910 12538
rect 14934 12486 14948 12538
rect 14948 12486 14960 12538
rect 14960 12486 14990 12538
rect 15014 12486 15024 12538
rect 15024 12486 15070 12538
rect 14774 12484 14830 12486
rect 14854 12484 14910 12486
rect 14934 12484 14990 12486
rect 15014 12484 15070 12486
rect 15290 13640 15346 13696
rect 14738 12144 14794 12200
rect 14922 12008 14978 12064
rect 14830 11872 14886 11928
rect 14774 11450 14830 11452
rect 14854 11450 14910 11452
rect 14934 11450 14990 11452
rect 15014 11450 15070 11452
rect 14774 11398 14820 11450
rect 14820 11398 14830 11450
rect 14854 11398 14884 11450
rect 14884 11398 14896 11450
rect 14896 11398 14910 11450
rect 14934 11398 14948 11450
rect 14948 11398 14960 11450
rect 14960 11398 14990 11450
rect 15014 11398 15024 11450
rect 15024 11398 15070 11450
rect 14774 11396 14830 11398
rect 14854 11396 14910 11398
rect 14934 11396 14990 11398
rect 15014 11396 15070 11398
rect 14922 11056 14978 11112
rect 14646 10920 14702 10976
rect 14830 10784 14886 10840
rect 15014 10648 15070 10704
rect 15382 13524 15438 13560
rect 15382 13504 15384 13524
rect 15384 13504 15436 13524
rect 15436 13504 15438 13524
rect 15382 13368 15438 13424
rect 15474 12824 15530 12880
rect 15382 12552 15438 12608
rect 15290 11192 15346 11248
rect 15198 10920 15254 10976
rect 14738 10512 14794 10568
rect 15290 10804 15346 10840
rect 15290 10784 15292 10804
rect 15292 10784 15344 10804
rect 15344 10784 15346 10804
rect 14774 10362 14830 10364
rect 14854 10362 14910 10364
rect 14934 10362 14990 10364
rect 15014 10362 15070 10364
rect 14774 10310 14820 10362
rect 14820 10310 14830 10362
rect 14854 10310 14884 10362
rect 14884 10310 14896 10362
rect 14896 10310 14910 10362
rect 14934 10310 14948 10362
rect 14948 10310 14960 10362
rect 14960 10310 14990 10362
rect 15014 10310 15024 10362
rect 15024 10310 15070 10362
rect 14774 10308 14830 10310
rect 14854 10308 14910 10310
rect 14934 10308 14990 10310
rect 15014 10308 15070 10310
rect 14554 9868 14556 9888
rect 14556 9868 14608 9888
rect 14608 9868 14610 9888
rect 14554 9832 14610 9868
rect 14830 9832 14886 9888
rect 14554 9288 14610 9344
rect 15106 9968 15162 10024
rect 15290 10240 15346 10296
rect 14554 9016 14610 9072
rect 14774 9274 14830 9276
rect 14854 9274 14910 9276
rect 14934 9274 14990 9276
rect 15014 9274 15070 9276
rect 14774 9222 14820 9274
rect 14820 9222 14830 9274
rect 14854 9222 14884 9274
rect 14884 9222 14896 9274
rect 14896 9222 14910 9274
rect 14934 9222 14948 9274
rect 14948 9222 14960 9274
rect 14960 9222 14990 9274
rect 15014 9222 15024 9274
rect 15024 9222 15070 9274
rect 14774 9220 14830 9222
rect 14854 9220 14910 9222
rect 14934 9220 14990 9222
rect 15014 9220 15070 9222
rect 14738 8744 14794 8800
rect 14738 8472 14794 8528
rect 14830 8336 14886 8392
rect 15106 8880 15162 8936
rect 15106 8356 15162 8392
rect 15106 8336 15108 8356
rect 15108 8336 15160 8356
rect 15160 8336 15162 8356
rect 14774 8186 14830 8188
rect 14854 8186 14910 8188
rect 14934 8186 14990 8188
rect 15014 8186 15070 8188
rect 14774 8134 14820 8186
rect 14820 8134 14830 8186
rect 14854 8134 14884 8186
rect 14884 8134 14896 8186
rect 14896 8134 14910 8186
rect 14934 8134 14948 8186
rect 14948 8134 14960 8186
rect 14960 8134 14990 8186
rect 15014 8134 15024 8186
rect 15024 8134 15070 8186
rect 14774 8132 14830 8134
rect 14854 8132 14910 8134
rect 14934 8132 14990 8134
rect 15014 8132 15070 8134
rect 14646 7792 14702 7848
rect 15106 7928 15162 7984
rect 14774 7098 14830 7100
rect 14854 7098 14910 7100
rect 14934 7098 14990 7100
rect 15014 7098 15070 7100
rect 14774 7046 14820 7098
rect 14820 7046 14830 7098
rect 14854 7046 14884 7098
rect 14884 7046 14896 7098
rect 14896 7046 14910 7098
rect 14934 7046 14948 7098
rect 14948 7046 14960 7098
rect 14960 7046 14990 7098
rect 15014 7046 15024 7098
rect 15024 7046 15070 7098
rect 14774 7044 14830 7046
rect 14854 7044 14910 7046
rect 14934 7044 14990 7046
rect 15014 7044 15070 7046
rect 14462 5752 14518 5808
rect 14462 5072 14518 5128
rect 14370 3848 14426 3904
rect 14774 6010 14830 6012
rect 14854 6010 14910 6012
rect 14934 6010 14990 6012
rect 15014 6010 15070 6012
rect 14774 5958 14820 6010
rect 14820 5958 14830 6010
rect 14854 5958 14884 6010
rect 14884 5958 14896 6010
rect 14896 5958 14910 6010
rect 14934 5958 14948 6010
rect 14948 5958 14960 6010
rect 14960 5958 14990 6010
rect 15014 5958 15024 6010
rect 15024 5958 15070 6010
rect 14774 5956 14830 5958
rect 14854 5956 14910 5958
rect 14934 5956 14990 5958
rect 15014 5956 15070 5958
rect 15658 13232 15714 13288
rect 15658 12144 15714 12200
rect 15474 10648 15530 10704
rect 15658 10376 15714 10432
rect 15566 10104 15622 10160
rect 15382 8880 15438 8936
rect 15198 5888 15254 5944
rect 15658 9696 15714 9752
rect 15566 6840 15622 6896
rect 15382 6296 15438 6352
rect 14774 4922 14830 4924
rect 14854 4922 14910 4924
rect 14934 4922 14990 4924
rect 15014 4922 15070 4924
rect 14774 4870 14820 4922
rect 14820 4870 14830 4922
rect 14854 4870 14884 4922
rect 14884 4870 14896 4922
rect 14896 4870 14910 4922
rect 14934 4870 14948 4922
rect 14948 4870 14960 4922
rect 14960 4870 14990 4922
rect 15014 4870 15024 4922
rect 15024 4870 15070 4922
rect 14774 4868 14830 4870
rect 14854 4868 14910 4870
rect 14934 4868 14990 4870
rect 15014 4868 15070 4870
rect 15290 5072 15346 5128
rect 14646 4392 14702 4448
rect 15014 3984 15070 4040
rect 14774 3834 14830 3836
rect 14854 3834 14910 3836
rect 14934 3834 14990 3836
rect 15014 3834 15070 3836
rect 14774 3782 14820 3834
rect 14820 3782 14830 3834
rect 14854 3782 14884 3834
rect 14884 3782 14896 3834
rect 14896 3782 14910 3834
rect 14934 3782 14948 3834
rect 14948 3782 14960 3834
rect 14960 3782 14990 3834
rect 15014 3782 15024 3834
rect 15024 3782 15070 3834
rect 14774 3780 14830 3782
rect 14854 3780 14910 3782
rect 14934 3780 14990 3782
rect 15014 3780 15070 3782
rect 14554 3440 14610 3496
rect 14774 2746 14830 2748
rect 14854 2746 14910 2748
rect 14934 2746 14990 2748
rect 15014 2746 15070 2748
rect 14774 2694 14820 2746
rect 14820 2694 14830 2746
rect 14854 2694 14884 2746
rect 14884 2694 14896 2746
rect 14896 2694 14910 2746
rect 14934 2694 14948 2746
rect 14948 2694 14960 2746
rect 14960 2694 14990 2746
rect 15014 2694 15024 2746
rect 15024 2694 15070 2746
rect 14774 2692 14830 2694
rect 14854 2692 14910 2694
rect 14934 2692 14990 2694
rect 15014 2692 15070 2694
rect 15290 2896 15346 2952
rect 14646 2352 14702 2408
rect 15014 2352 15070 2408
rect 14830 2080 14886 2136
rect 14554 1944 14610 2000
rect 15750 8372 15752 8392
rect 15752 8372 15804 8392
rect 15804 8372 15806 8392
rect 15750 8336 15806 8372
rect 15750 5208 15806 5264
rect 15658 3168 15714 3224
rect 15750 3032 15806 3088
rect 16026 4140 16082 4176
rect 16026 4120 16028 4140
rect 16028 4120 16080 4140
rect 16080 4120 16082 4140
rect 16394 9424 16450 9480
rect 16302 7384 16358 7440
rect 16302 6840 16358 6896
rect 16026 2488 16082 2544
rect 14774 1658 14830 1660
rect 14854 1658 14910 1660
rect 14934 1658 14990 1660
rect 15014 1658 15070 1660
rect 14774 1606 14820 1658
rect 14820 1606 14830 1658
rect 14854 1606 14884 1658
rect 14884 1606 14896 1658
rect 14896 1606 14910 1658
rect 14934 1606 14948 1658
rect 14948 1606 14960 1658
rect 14960 1606 14990 1658
rect 15014 1606 15024 1658
rect 15024 1606 15070 1658
rect 14774 1604 14830 1606
rect 14854 1604 14910 1606
rect 14934 1604 14990 1606
rect 15014 1604 15070 1606
rect 14370 1400 14426 1456
rect 14186 856 14242 912
rect 14094 720 14150 776
rect 17222 4256 17278 4312
rect 17498 13096 17554 13152
rect 17682 6704 17738 6760
rect 17590 3304 17646 3360
<< metal3 >>
rect 0 23218 400 23248
rect 1577 23218 1643 23221
rect 0 23216 1643 23218
rect 0 23160 1582 23216
rect 1638 23160 1643 23216
rect 0 23158 1643 23160
rect 0 23128 400 23158
rect 1577 23155 1643 23158
rect 4894 22880 5210 22881
rect 4894 22816 4900 22880
rect 4964 22816 4980 22880
rect 5044 22816 5060 22880
rect 5124 22816 5140 22880
rect 5204 22816 5210 22880
rect 4894 22815 5210 22816
rect 8842 22880 9158 22881
rect 8842 22816 8848 22880
rect 8912 22816 8928 22880
rect 8992 22816 9008 22880
rect 9072 22816 9088 22880
rect 9152 22816 9158 22880
rect 8842 22815 9158 22816
rect 12790 22880 13106 22881
rect 12790 22816 12796 22880
rect 12860 22816 12876 22880
rect 12940 22816 12956 22880
rect 13020 22816 13036 22880
rect 13100 22816 13106 22880
rect 12790 22815 13106 22816
rect 1485 22538 1551 22541
rect 16614 22538 16620 22540
rect 1485 22536 16620 22538
rect 1485 22480 1490 22536
rect 1546 22480 16620 22536
rect 1485 22478 16620 22480
rect 1485 22475 1551 22478
rect 16614 22476 16620 22478
rect 16684 22476 16690 22540
rect 2920 22336 3236 22337
rect 2920 22272 2926 22336
rect 2990 22272 3006 22336
rect 3070 22272 3086 22336
rect 3150 22272 3166 22336
rect 3230 22272 3236 22336
rect 2920 22271 3236 22272
rect 6868 22336 7184 22337
rect 6868 22272 6874 22336
rect 6938 22272 6954 22336
rect 7018 22272 7034 22336
rect 7098 22272 7114 22336
rect 7178 22272 7184 22336
rect 6868 22271 7184 22272
rect 10816 22336 11132 22337
rect 10816 22272 10822 22336
rect 10886 22272 10902 22336
rect 10966 22272 10982 22336
rect 11046 22272 11062 22336
rect 11126 22272 11132 22336
rect 10816 22271 11132 22272
rect 14764 22336 15080 22337
rect 14764 22272 14770 22336
rect 14834 22272 14850 22336
rect 14914 22272 14930 22336
rect 14994 22272 15010 22336
rect 15074 22272 15080 22336
rect 14764 22271 15080 22272
rect 4894 21792 5210 21793
rect 0 21722 400 21752
rect 4894 21728 4900 21792
rect 4964 21728 4980 21792
rect 5044 21728 5060 21792
rect 5124 21728 5140 21792
rect 5204 21728 5210 21792
rect 4894 21727 5210 21728
rect 8842 21792 9158 21793
rect 8842 21728 8848 21792
rect 8912 21728 8928 21792
rect 8992 21728 9008 21792
rect 9072 21728 9088 21792
rect 9152 21728 9158 21792
rect 8842 21727 9158 21728
rect 12790 21792 13106 21793
rect 12790 21728 12796 21792
rect 12860 21728 12876 21792
rect 12940 21728 12956 21792
rect 13020 21728 13036 21792
rect 13100 21728 13106 21792
rect 12790 21727 13106 21728
rect 2405 21722 2471 21725
rect 0 21720 2471 21722
rect 0 21664 2410 21720
rect 2466 21664 2471 21720
rect 0 21662 2471 21664
rect 0 21632 400 21662
rect 2405 21659 2471 21662
rect 2920 21248 3236 21249
rect 2920 21184 2926 21248
rect 2990 21184 3006 21248
rect 3070 21184 3086 21248
rect 3150 21184 3166 21248
rect 3230 21184 3236 21248
rect 2920 21183 3236 21184
rect 6868 21248 7184 21249
rect 6868 21184 6874 21248
rect 6938 21184 6954 21248
rect 7018 21184 7034 21248
rect 7098 21184 7114 21248
rect 7178 21184 7184 21248
rect 6868 21183 7184 21184
rect 10816 21248 11132 21249
rect 10816 21184 10822 21248
rect 10886 21184 10902 21248
rect 10966 21184 10982 21248
rect 11046 21184 11062 21248
rect 11126 21184 11132 21248
rect 10816 21183 11132 21184
rect 14764 21248 15080 21249
rect 14764 21184 14770 21248
rect 14834 21184 14850 21248
rect 14914 21184 14930 21248
rect 14994 21184 15010 21248
rect 15074 21184 15080 21248
rect 14764 21183 15080 21184
rect 4894 20704 5210 20705
rect 4894 20640 4900 20704
rect 4964 20640 4980 20704
rect 5044 20640 5060 20704
rect 5124 20640 5140 20704
rect 5204 20640 5210 20704
rect 4894 20639 5210 20640
rect 8842 20704 9158 20705
rect 8842 20640 8848 20704
rect 8912 20640 8928 20704
rect 8992 20640 9008 20704
rect 9072 20640 9088 20704
rect 9152 20640 9158 20704
rect 8842 20639 9158 20640
rect 12790 20704 13106 20705
rect 12790 20640 12796 20704
rect 12860 20640 12876 20704
rect 12940 20640 12956 20704
rect 13020 20640 13036 20704
rect 13100 20640 13106 20704
rect 12790 20639 13106 20640
rect 3141 20362 3207 20365
rect 3734 20362 3740 20364
rect 3141 20360 3740 20362
rect 3141 20304 3146 20360
rect 3202 20304 3740 20360
rect 3141 20302 3740 20304
rect 3141 20299 3207 20302
rect 3734 20300 3740 20302
rect 3804 20362 3810 20364
rect 4337 20362 4403 20365
rect 3804 20360 4403 20362
rect 3804 20304 4342 20360
rect 4398 20304 4403 20360
rect 3804 20302 4403 20304
rect 3804 20300 3810 20302
rect 4337 20299 4403 20302
rect 0 20226 400 20256
rect 2773 20226 2839 20229
rect 0 20224 2839 20226
rect 0 20168 2778 20224
rect 2834 20168 2839 20224
rect 0 20166 2839 20168
rect 0 20136 400 20166
rect 2773 20163 2839 20166
rect 3601 20226 3667 20229
rect 5809 20226 5875 20229
rect 3601 20224 5875 20226
rect 3601 20168 3606 20224
rect 3662 20168 5814 20224
rect 5870 20168 5875 20224
rect 3601 20166 5875 20168
rect 3601 20163 3667 20166
rect 5809 20163 5875 20166
rect 2920 20160 3236 20161
rect 2920 20096 2926 20160
rect 2990 20096 3006 20160
rect 3070 20096 3086 20160
rect 3150 20096 3166 20160
rect 3230 20096 3236 20160
rect 2920 20095 3236 20096
rect 6868 20160 7184 20161
rect 6868 20096 6874 20160
rect 6938 20096 6954 20160
rect 7018 20096 7034 20160
rect 7098 20096 7114 20160
rect 7178 20096 7184 20160
rect 6868 20095 7184 20096
rect 10816 20160 11132 20161
rect 10816 20096 10822 20160
rect 10886 20096 10902 20160
rect 10966 20096 10982 20160
rect 11046 20096 11062 20160
rect 11126 20096 11132 20160
rect 10816 20095 11132 20096
rect 14764 20160 15080 20161
rect 14764 20096 14770 20160
rect 14834 20096 14850 20160
rect 14914 20096 14930 20160
rect 14994 20096 15010 20160
rect 15074 20096 15080 20160
rect 14764 20095 15080 20096
rect 3785 20090 3851 20093
rect 3328 20088 3851 20090
rect 3328 20032 3790 20088
rect 3846 20032 3851 20088
rect 3328 20030 3851 20032
rect 3141 19954 3207 19957
rect 3328 19954 3388 20030
rect 3785 20027 3851 20030
rect 4705 20090 4771 20093
rect 5533 20090 5599 20093
rect 4705 20088 5599 20090
rect 4705 20032 4710 20088
rect 4766 20032 5538 20088
rect 5594 20032 5599 20088
rect 4705 20030 5599 20032
rect 4705 20027 4771 20030
rect 5533 20027 5599 20030
rect 3141 19952 3388 19954
rect 3141 19896 3146 19952
rect 3202 19896 3388 19952
rect 3141 19894 3388 19896
rect 3969 19954 4035 19957
rect 6085 19954 6151 19957
rect 3969 19952 6151 19954
rect 3969 19896 3974 19952
rect 4030 19896 6090 19952
rect 6146 19896 6151 19952
rect 3969 19894 6151 19896
rect 3141 19891 3207 19894
rect 3969 19891 4035 19894
rect 6085 19891 6151 19894
rect 2865 19818 2931 19821
rect 5441 19818 5507 19821
rect 6637 19818 6703 19821
rect 2865 19816 6703 19818
rect 2865 19760 2870 19816
rect 2926 19760 5446 19816
rect 5502 19760 6642 19816
rect 6698 19760 6703 19816
rect 2865 19758 6703 19760
rect 2865 19755 2931 19758
rect 5441 19755 5507 19758
rect 6637 19755 6703 19758
rect 3325 19682 3391 19685
rect 4705 19682 4771 19685
rect 3325 19680 4771 19682
rect 3325 19624 3330 19680
rect 3386 19624 4710 19680
rect 4766 19624 4771 19680
rect 3325 19622 4771 19624
rect 3325 19619 3391 19622
rect 4705 19619 4771 19622
rect 5625 19682 5691 19685
rect 8661 19682 8727 19685
rect 5625 19680 8727 19682
rect 5625 19624 5630 19680
rect 5686 19624 8666 19680
rect 8722 19624 8727 19680
rect 5625 19622 8727 19624
rect 5625 19619 5691 19622
rect 8661 19619 8727 19622
rect 4894 19616 5210 19617
rect 4894 19552 4900 19616
rect 4964 19552 4980 19616
rect 5044 19552 5060 19616
rect 5124 19552 5140 19616
rect 5204 19552 5210 19616
rect 4894 19551 5210 19552
rect 8842 19616 9158 19617
rect 8842 19552 8848 19616
rect 8912 19552 8928 19616
rect 8992 19552 9008 19616
rect 9072 19552 9088 19616
rect 9152 19552 9158 19616
rect 8842 19551 9158 19552
rect 12790 19616 13106 19617
rect 12790 19552 12796 19616
rect 12860 19552 12876 19616
rect 12940 19552 12956 19616
rect 13020 19552 13036 19616
rect 13100 19552 13106 19616
rect 12790 19551 13106 19552
rect 5901 19546 5967 19549
rect 5901 19544 8770 19546
rect 5901 19488 5906 19544
rect 5962 19488 8770 19544
rect 5901 19486 8770 19488
rect 5901 19483 5967 19486
rect 2589 19410 2655 19413
rect 4705 19410 4771 19413
rect 2589 19408 4771 19410
rect 2589 19352 2594 19408
rect 2650 19352 4710 19408
rect 4766 19352 4771 19408
rect 2589 19350 4771 19352
rect 2589 19347 2655 19350
rect 4705 19347 4771 19350
rect 5257 19410 5323 19413
rect 6545 19410 6611 19413
rect 5257 19408 6611 19410
rect 5257 19352 5262 19408
rect 5318 19352 6550 19408
rect 6606 19352 6611 19408
rect 5257 19350 6611 19352
rect 8710 19410 8770 19486
rect 9213 19410 9279 19413
rect 8710 19408 9279 19410
rect 8710 19352 9218 19408
rect 9274 19352 9279 19408
rect 8710 19350 9279 19352
rect 5257 19347 5323 19350
rect 6545 19347 6611 19350
rect 9213 19347 9279 19350
rect 473 19274 539 19277
rect 3325 19274 3391 19277
rect 473 19272 3391 19274
rect 473 19216 478 19272
rect 534 19216 3330 19272
rect 3386 19216 3391 19272
rect 473 19214 3391 19216
rect 473 19211 539 19214
rect 3325 19211 3391 19214
rect 4470 19212 4476 19276
rect 4540 19274 4546 19276
rect 4705 19274 4771 19277
rect 4540 19272 4771 19274
rect 4540 19216 4710 19272
rect 4766 19216 4771 19272
rect 4540 19214 4771 19216
rect 4540 19212 4546 19214
rect 4705 19211 4771 19214
rect 2920 19072 3236 19073
rect 2920 19008 2926 19072
rect 2990 19008 3006 19072
rect 3070 19008 3086 19072
rect 3150 19008 3166 19072
rect 3230 19008 3236 19072
rect 2920 19007 3236 19008
rect 6868 19072 7184 19073
rect 6868 19008 6874 19072
rect 6938 19008 6954 19072
rect 7018 19008 7034 19072
rect 7098 19008 7114 19072
rect 7178 19008 7184 19072
rect 6868 19007 7184 19008
rect 10816 19072 11132 19073
rect 10816 19008 10822 19072
rect 10886 19008 10902 19072
rect 10966 19008 10982 19072
rect 11046 19008 11062 19072
rect 11126 19008 11132 19072
rect 10816 19007 11132 19008
rect 14764 19072 15080 19073
rect 14764 19008 14770 19072
rect 14834 19008 14850 19072
rect 14914 19008 14930 19072
rect 14994 19008 15010 19072
rect 15074 19008 15080 19072
rect 14764 19007 15080 19008
rect 6085 19002 6151 19005
rect 3328 19000 6151 19002
rect 3328 18944 6090 19000
rect 6146 18944 6151 19000
rect 3328 18942 6151 18944
rect 2589 18866 2655 18869
rect 3328 18866 3388 18942
rect 6085 18939 6151 18942
rect 2589 18864 3388 18866
rect 2589 18808 2594 18864
rect 2650 18808 3388 18864
rect 2589 18806 3388 18808
rect 4061 18866 4127 18869
rect 4654 18866 4660 18868
rect 4061 18864 4660 18866
rect 4061 18808 4066 18864
rect 4122 18808 4660 18864
rect 4061 18806 4660 18808
rect 2589 18803 2655 18806
rect 4061 18803 4127 18806
rect 4654 18804 4660 18806
rect 4724 18804 4730 18868
rect 5717 18866 5783 18869
rect 8477 18866 8543 18869
rect 5717 18864 8543 18866
rect 5717 18808 5722 18864
rect 5778 18808 8482 18864
rect 8538 18808 8543 18864
rect 5717 18806 8543 18808
rect 5717 18803 5783 18806
rect 8477 18803 8543 18806
rect 0 18730 400 18760
rect 3693 18730 3759 18733
rect 0 18728 3759 18730
rect 0 18672 3698 18728
rect 3754 18672 3759 18728
rect 0 18670 3759 18672
rect 0 18640 400 18670
rect 3693 18667 3759 18670
rect 5758 18668 5764 18732
rect 5828 18730 5834 18732
rect 8477 18730 8543 18733
rect 15193 18730 15259 18733
rect 5828 18728 8543 18730
rect 5828 18672 8482 18728
rect 8538 18672 8543 18728
rect 5828 18670 8543 18672
rect 5828 18668 5834 18670
rect 8477 18667 8543 18670
rect 8664 18728 15259 18730
rect 8664 18672 15198 18728
rect 15254 18672 15259 18728
rect 8664 18670 15259 18672
rect 2446 18532 2452 18596
rect 2516 18594 2522 18596
rect 3049 18594 3115 18597
rect 2516 18592 3115 18594
rect 2516 18536 3054 18592
rect 3110 18536 3115 18592
rect 2516 18534 3115 18536
rect 2516 18532 2522 18534
rect 3049 18531 3115 18534
rect 7649 18594 7715 18597
rect 8664 18594 8724 18670
rect 15193 18667 15259 18670
rect 12065 18594 12131 18597
rect 7649 18592 8724 18594
rect 7649 18536 7654 18592
rect 7710 18536 8724 18592
rect 7649 18534 8724 18536
rect 9308 18592 12131 18594
rect 9308 18536 12070 18592
rect 12126 18536 12131 18592
rect 9308 18534 12131 18536
rect 7649 18531 7715 18534
rect 4894 18528 5210 18529
rect 4894 18464 4900 18528
rect 4964 18464 4980 18528
rect 5044 18464 5060 18528
rect 5124 18464 5140 18528
rect 5204 18464 5210 18528
rect 4894 18463 5210 18464
rect 8842 18528 9158 18529
rect 8842 18464 8848 18528
rect 8912 18464 8928 18528
rect 8992 18464 9008 18528
rect 9072 18464 9088 18528
rect 9152 18464 9158 18528
rect 8842 18463 9158 18464
rect 3785 18458 3851 18461
rect 4705 18458 4771 18461
rect 8702 18458 8708 18460
rect 3785 18456 4771 18458
rect 3785 18400 3790 18456
rect 3846 18400 4710 18456
rect 4766 18400 4771 18456
rect 3785 18398 4771 18400
rect 3785 18395 3851 18398
rect 4705 18395 4771 18398
rect 5398 18398 8708 18458
rect 1710 18260 1716 18324
rect 1780 18322 1786 18324
rect 5398 18322 5458 18398
rect 8702 18396 8708 18398
rect 8772 18396 8778 18460
rect 1780 18262 5458 18322
rect 1780 18260 1786 18262
rect 5942 18260 5948 18324
rect 6012 18322 6018 18324
rect 6269 18322 6335 18325
rect 6012 18320 6335 18322
rect 6012 18264 6274 18320
rect 6330 18264 6335 18320
rect 6012 18262 6335 18264
rect 6012 18260 6018 18262
rect 6269 18259 6335 18262
rect 7097 18322 7163 18325
rect 7782 18322 7788 18324
rect 7097 18320 7788 18322
rect 7097 18264 7102 18320
rect 7158 18264 7788 18320
rect 7097 18262 7788 18264
rect 7097 18259 7163 18262
rect 7782 18260 7788 18262
rect 7852 18260 7858 18324
rect 7925 18322 7991 18325
rect 9308 18322 9368 18534
rect 12065 18531 12131 18534
rect 12790 18528 13106 18529
rect 12790 18464 12796 18528
rect 12860 18464 12876 18528
rect 12940 18464 12956 18528
rect 13020 18464 13036 18528
rect 13100 18464 13106 18528
rect 12790 18463 13106 18464
rect 10777 18458 10843 18461
rect 11462 18458 11468 18460
rect 10777 18456 11468 18458
rect 10777 18400 10782 18456
rect 10838 18400 11468 18456
rect 10777 18398 11468 18400
rect 10777 18395 10843 18398
rect 11462 18396 11468 18398
rect 11532 18396 11538 18460
rect 7925 18320 9368 18322
rect 7925 18264 7930 18320
rect 7986 18264 9368 18320
rect 7925 18262 9368 18264
rect 9489 18322 9555 18325
rect 16798 18322 16804 18324
rect 9489 18320 16804 18322
rect 9489 18264 9494 18320
rect 9550 18264 16804 18320
rect 9489 18262 16804 18264
rect 7925 18259 7991 18262
rect 9489 18259 9555 18262
rect 16798 18260 16804 18262
rect 16868 18260 16874 18324
rect 2681 18186 2747 18189
rect 4061 18186 4127 18189
rect 5625 18186 5691 18189
rect 12566 18186 12572 18188
rect 2681 18184 4538 18186
rect 2681 18128 2686 18184
rect 2742 18128 4066 18184
rect 4122 18128 4538 18184
rect 2681 18126 4538 18128
rect 2681 18123 2747 18126
rect 4061 18123 4127 18126
rect 4061 18052 4127 18053
rect 4061 18048 4108 18052
rect 4172 18050 4178 18052
rect 4061 17992 4066 18048
rect 4061 17988 4108 17992
rect 4172 17990 4218 18050
rect 4172 17988 4178 17990
rect 4061 17987 4127 17988
rect 2920 17984 3236 17985
rect 2920 17920 2926 17984
rect 2990 17920 3006 17984
rect 3070 17920 3086 17984
rect 3150 17920 3166 17984
rect 3230 17920 3236 17984
rect 2920 17919 3236 17920
rect 4478 17914 4538 18126
rect 5625 18184 12572 18186
rect 5625 18128 5630 18184
rect 5686 18128 12572 18184
rect 5625 18126 12572 18128
rect 5625 18123 5691 18126
rect 12566 18124 12572 18126
rect 12636 18124 12642 18188
rect 6126 17988 6132 18052
rect 6196 18050 6202 18052
rect 6545 18050 6611 18053
rect 6196 18048 6611 18050
rect 6196 17992 6550 18048
rect 6606 17992 6611 18048
rect 6196 17990 6611 17992
rect 6196 17988 6202 17990
rect 6545 17987 6611 17990
rect 8109 18050 8175 18053
rect 9254 18050 9260 18052
rect 8109 18048 9260 18050
rect 8109 17992 8114 18048
rect 8170 17992 9260 18048
rect 8109 17990 9260 17992
rect 8109 17987 8175 17990
rect 9254 17988 9260 17990
rect 9324 17988 9330 18052
rect 9673 18050 9739 18053
rect 9806 18050 9812 18052
rect 9673 18048 9812 18050
rect 9673 17992 9678 18048
rect 9734 17992 9812 18048
rect 9673 17990 9812 17992
rect 9673 17987 9739 17990
rect 9806 17988 9812 17990
rect 9876 17988 9882 18052
rect 6868 17984 7184 17985
rect 6868 17920 6874 17984
rect 6938 17920 6954 17984
rect 7018 17920 7034 17984
rect 7098 17920 7114 17984
rect 7178 17920 7184 17984
rect 6868 17919 7184 17920
rect 10816 17984 11132 17985
rect 10816 17920 10822 17984
rect 10886 17920 10902 17984
rect 10966 17920 10982 17984
rect 11046 17920 11062 17984
rect 11126 17920 11132 17984
rect 10816 17919 11132 17920
rect 14764 17984 15080 17985
rect 14764 17920 14770 17984
rect 14834 17920 14850 17984
rect 14914 17920 14930 17984
rect 14994 17920 15010 17984
rect 15074 17920 15080 17984
rect 14764 17919 15080 17920
rect 6361 17914 6427 17917
rect 4478 17912 6427 17914
rect 4478 17856 6366 17912
rect 6422 17856 6427 17912
rect 4478 17854 6427 17856
rect 6361 17851 6427 17854
rect 7925 17914 7991 17917
rect 8150 17914 8156 17916
rect 7925 17912 8156 17914
rect 7925 17856 7930 17912
rect 7986 17856 8156 17912
rect 7925 17854 8156 17856
rect 7925 17851 7991 17854
rect 8150 17852 8156 17854
rect 8220 17914 8226 17916
rect 8220 17854 9690 17914
rect 8220 17852 8226 17854
rect 13 17778 79 17781
rect 9397 17778 9463 17781
rect 13 17776 9463 17778
rect 13 17720 18 17776
rect 74 17720 9402 17776
rect 9458 17720 9463 17776
rect 13 17718 9463 17720
rect 9630 17778 9690 17854
rect 11513 17778 11579 17781
rect 9630 17776 11579 17778
rect 9630 17720 11518 17776
rect 11574 17720 11579 17776
rect 9630 17718 11579 17720
rect 13 17715 79 17718
rect 9397 17715 9463 17718
rect 11513 17715 11579 17718
rect 933 17642 999 17645
rect 5165 17642 5231 17645
rect 933 17640 5231 17642
rect 933 17584 938 17640
rect 994 17584 5170 17640
rect 5226 17584 5231 17640
rect 933 17582 5231 17584
rect 933 17579 999 17582
rect 5165 17579 5231 17582
rect 7097 17642 7163 17645
rect 11145 17642 11211 17645
rect 7097 17640 11211 17642
rect 7097 17584 7102 17640
rect 7158 17584 11150 17640
rect 11206 17584 11211 17640
rect 7097 17582 11211 17584
rect 7097 17579 7163 17582
rect 11145 17579 11211 17582
rect 6361 17506 6427 17509
rect 7649 17506 7715 17509
rect 6361 17504 7715 17506
rect 6361 17448 6366 17504
rect 6422 17448 7654 17504
rect 7710 17448 7715 17504
rect 6361 17446 7715 17448
rect 6361 17443 6427 17446
rect 7649 17443 7715 17446
rect 8201 17506 8267 17509
rect 8569 17506 8635 17509
rect 8201 17504 8635 17506
rect 8201 17448 8206 17504
rect 8262 17448 8574 17504
rect 8630 17448 8635 17504
rect 8201 17446 8635 17448
rect 8201 17443 8267 17446
rect 8569 17443 8635 17446
rect 9857 17506 9923 17509
rect 11646 17506 11652 17508
rect 9857 17504 11652 17506
rect 9857 17448 9862 17504
rect 9918 17448 11652 17504
rect 9857 17446 11652 17448
rect 9857 17443 9923 17446
rect 11646 17444 11652 17446
rect 11716 17444 11722 17508
rect 4894 17440 5210 17441
rect 4894 17376 4900 17440
rect 4964 17376 4980 17440
rect 5044 17376 5060 17440
rect 5124 17376 5140 17440
rect 5204 17376 5210 17440
rect 4894 17375 5210 17376
rect 8842 17440 9158 17441
rect 8842 17376 8848 17440
rect 8912 17376 8928 17440
rect 8992 17376 9008 17440
rect 9072 17376 9088 17440
rect 9152 17376 9158 17440
rect 8842 17375 9158 17376
rect 12790 17440 13106 17441
rect 12790 17376 12796 17440
rect 12860 17376 12876 17440
rect 12940 17376 12956 17440
rect 13020 17376 13036 17440
rect 13100 17376 13106 17440
rect 12790 17375 13106 17376
rect 7373 17370 7439 17373
rect 8293 17370 8359 17373
rect 7373 17368 8359 17370
rect 7373 17312 7378 17368
rect 7434 17312 8298 17368
rect 8354 17312 8359 17368
rect 7373 17310 8359 17312
rect 7373 17307 7439 17310
rect 8293 17307 8359 17310
rect 10041 17370 10107 17373
rect 10542 17370 10548 17372
rect 10041 17368 10548 17370
rect 10041 17312 10046 17368
rect 10102 17312 10548 17368
rect 10041 17310 10548 17312
rect 10041 17307 10107 17310
rect 10542 17308 10548 17310
rect 10612 17308 10618 17372
rect 0 17234 400 17264
rect 3325 17234 3391 17237
rect 0 17232 3391 17234
rect 0 17176 3330 17232
rect 3386 17176 3391 17232
rect 0 17174 3391 17176
rect 0 17144 400 17174
rect 3325 17171 3391 17174
rect 3918 17172 3924 17236
rect 3988 17234 3994 17236
rect 4337 17234 4403 17237
rect 3988 17232 4403 17234
rect 3988 17176 4342 17232
rect 4398 17176 4403 17232
rect 3988 17174 4403 17176
rect 3988 17172 3994 17174
rect 4337 17171 4403 17174
rect 6453 17234 6519 17237
rect 12341 17234 12407 17237
rect 6453 17232 12407 17234
rect 6453 17176 6458 17232
rect 6514 17176 12346 17232
rect 12402 17176 12407 17232
rect 6453 17174 12407 17176
rect 6453 17171 6519 17174
rect 12341 17171 12407 17174
rect 6494 17036 6500 17100
rect 6564 17098 6570 17100
rect 9029 17098 9095 17101
rect 6564 17096 9095 17098
rect 6564 17040 9034 17096
rect 9090 17040 9095 17096
rect 6564 17038 9095 17040
rect 6564 17036 6570 17038
rect 9029 17035 9095 17038
rect 9438 17036 9444 17100
rect 9508 17098 9514 17100
rect 9673 17098 9739 17101
rect 9806 17098 9812 17100
rect 9508 17096 9812 17098
rect 9508 17040 9678 17096
rect 9734 17040 9812 17096
rect 9508 17038 9812 17040
rect 9508 17036 9514 17038
rect 9673 17035 9739 17038
rect 9806 17036 9812 17038
rect 9876 17036 9882 17100
rect 10041 17098 10107 17101
rect 14038 17098 14044 17100
rect 10041 17096 14044 17098
rect 10041 17040 10046 17096
rect 10102 17040 14044 17096
rect 10041 17038 14044 17040
rect 10041 17035 10107 17038
rect 14038 17036 14044 17038
rect 14108 17036 14114 17100
rect 7966 16900 7972 16964
rect 8036 16962 8042 16964
rect 8477 16962 8543 16965
rect 9489 16962 9555 16965
rect 8036 16960 9555 16962
rect 8036 16904 8482 16960
rect 8538 16904 9494 16960
rect 9550 16904 9555 16960
rect 8036 16902 9555 16904
rect 8036 16900 8042 16902
rect 8477 16899 8543 16902
rect 9489 16899 9555 16902
rect 9673 16962 9739 16965
rect 10685 16962 10751 16965
rect 9673 16960 10751 16962
rect 9673 16904 9678 16960
rect 9734 16904 10690 16960
rect 10746 16904 10751 16960
rect 9673 16902 10751 16904
rect 9673 16899 9739 16902
rect 10685 16899 10751 16902
rect 2920 16896 3236 16897
rect 2920 16832 2926 16896
rect 2990 16832 3006 16896
rect 3070 16832 3086 16896
rect 3150 16832 3166 16896
rect 3230 16832 3236 16896
rect 2920 16831 3236 16832
rect 6868 16896 7184 16897
rect 6868 16832 6874 16896
rect 6938 16832 6954 16896
rect 7018 16832 7034 16896
rect 7098 16832 7114 16896
rect 7178 16832 7184 16896
rect 6868 16831 7184 16832
rect 10816 16896 11132 16897
rect 10816 16832 10822 16896
rect 10886 16832 10902 16896
rect 10966 16832 10982 16896
rect 11046 16832 11062 16896
rect 11126 16832 11132 16896
rect 10816 16831 11132 16832
rect 14764 16896 15080 16897
rect 14764 16832 14770 16896
rect 14834 16832 14850 16896
rect 14914 16832 14930 16896
rect 14994 16832 15010 16896
rect 15074 16832 15080 16896
rect 14764 16831 15080 16832
rect 5441 16828 5507 16829
rect 5390 16826 5396 16828
rect 5350 16766 5396 16826
rect 5460 16824 5507 16828
rect 5502 16768 5507 16824
rect 5390 16764 5396 16766
rect 5460 16764 5507 16768
rect 5441 16763 5507 16764
rect 7465 16826 7531 16829
rect 7925 16826 7991 16829
rect 7465 16824 7991 16826
rect 7465 16768 7470 16824
rect 7526 16768 7930 16824
rect 7986 16768 7991 16824
rect 7465 16766 7991 16768
rect 7465 16763 7531 16766
rect 7925 16763 7991 16766
rect 8702 16764 8708 16828
rect 8772 16826 8778 16828
rect 10593 16826 10659 16829
rect 8772 16824 10659 16826
rect 8772 16768 10598 16824
rect 10654 16768 10659 16824
rect 8772 16766 10659 16768
rect 8772 16764 8778 16766
rect 10593 16763 10659 16766
rect 2446 16628 2452 16692
rect 2516 16690 2522 16692
rect 6913 16690 6979 16693
rect 2516 16688 6979 16690
rect 2516 16632 6918 16688
rect 6974 16632 6979 16688
rect 2516 16630 6979 16632
rect 2516 16628 2522 16630
rect 6913 16627 6979 16630
rect 7598 16628 7604 16692
rect 7668 16690 7674 16692
rect 7833 16690 7899 16693
rect 7668 16688 7899 16690
rect 7668 16632 7838 16688
rect 7894 16632 7899 16688
rect 7668 16630 7899 16632
rect 7668 16628 7674 16630
rect 7833 16627 7899 16630
rect 8518 16628 8524 16692
rect 8588 16690 8594 16692
rect 11697 16690 11763 16693
rect 8588 16688 11763 16690
rect 8588 16632 11702 16688
rect 11758 16632 11763 16688
rect 8588 16630 11763 16632
rect 8588 16628 8594 16630
rect 11697 16627 11763 16630
rect 2262 16492 2268 16556
rect 2332 16554 2338 16556
rect 2405 16554 2471 16557
rect 2332 16552 2471 16554
rect 2332 16496 2410 16552
rect 2466 16496 2471 16552
rect 2332 16494 2471 16496
rect 2332 16492 2338 16494
rect 2405 16491 2471 16494
rect 2681 16554 2747 16557
rect 3366 16554 3372 16556
rect 2681 16552 3372 16554
rect 2681 16496 2686 16552
rect 2742 16496 3372 16552
rect 2681 16494 3372 16496
rect 2681 16491 2747 16494
rect 3366 16492 3372 16494
rect 3436 16492 3442 16556
rect 4797 16554 4863 16557
rect 7373 16556 7439 16557
rect 5574 16554 5580 16556
rect 4797 16552 5580 16554
rect 4797 16496 4802 16552
rect 4858 16496 5580 16552
rect 4797 16494 5580 16496
rect 4797 16491 4863 16494
rect 5574 16492 5580 16494
rect 5644 16492 5650 16556
rect 7373 16552 7420 16556
rect 7484 16554 7490 16556
rect 8293 16554 8359 16557
rect 10593 16554 10659 16557
rect 7373 16496 7378 16552
rect 7373 16492 7420 16496
rect 7484 16494 7530 16554
rect 7606 16552 10659 16554
rect 7606 16496 8298 16552
rect 8354 16496 10598 16552
rect 10654 16496 10659 16552
rect 7606 16494 10659 16496
rect 7484 16492 7490 16494
rect 7373 16491 7439 16492
rect 1945 16418 2011 16421
rect 2405 16418 2471 16421
rect 1945 16416 2471 16418
rect 1945 16360 1950 16416
rect 2006 16360 2410 16416
rect 2466 16360 2471 16416
rect 1945 16358 2471 16360
rect 1945 16355 2011 16358
rect 2405 16355 2471 16358
rect 2630 16356 2636 16420
rect 2700 16418 2706 16420
rect 4521 16418 4587 16421
rect 6729 16420 6795 16421
rect 2700 16416 4587 16418
rect 2700 16360 4526 16416
rect 4582 16360 4587 16416
rect 2700 16358 4587 16360
rect 2700 16356 2706 16358
rect 4521 16355 4587 16358
rect 6678 16356 6684 16420
rect 6748 16418 6795 16420
rect 6748 16416 6840 16418
rect 6790 16360 6840 16416
rect 6748 16358 6840 16360
rect 6748 16356 6795 16358
rect 6729 16355 6795 16356
rect 4894 16352 5210 16353
rect 4894 16288 4900 16352
rect 4964 16288 4980 16352
rect 5044 16288 5060 16352
rect 5124 16288 5140 16352
rect 5204 16288 5210 16352
rect 4894 16287 5210 16288
rect 565 16282 631 16285
rect 565 16280 4400 16282
rect 565 16224 570 16280
rect 626 16224 4400 16280
rect 565 16222 4400 16224
rect 565 16219 631 16222
rect 4340 16146 4400 16222
rect 6310 16220 6316 16284
rect 6380 16282 6386 16284
rect 6637 16282 6703 16285
rect 6380 16280 6703 16282
rect 6380 16224 6642 16280
rect 6698 16224 6703 16280
rect 6380 16222 6703 16224
rect 6380 16220 6386 16222
rect 6637 16219 6703 16222
rect 7281 16282 7347 16285
rect 7606 16282 7666 16494
rect 8293 16491 8359 16494
rect 10593 16491 10659 16494
rect 9673 16418 9739 16421
rect 9949 16420 10015 16421
rect 9806 16418 9812 16420
rect 9673 16416 9812 16418
rect 9673 16360 9678 16416
rect 9734 16360 9812 16416
rect 9673 16358 9812 16360
rect 9673 16355 9739 16358
rect 9806 16356 9812 16358
rect 9876 16356 9882 16420
rect 9949 16416 9996 16420
rect 10060 16418 10066 16420
rect 10501 16418 10567 16421
rect 12014 16418 12020 16420
rect 9949 16360 9954 16416
rect 9949 16356 9996 16360
rect 10060 16358 10106 16418
rect 10501 16416 12020 16418
rect 10501 16360 10506 16416
rect 10562 16360 12020 16416
rect 10501 16358 12020 16360
rect 10060 16356 10066 16358
rect 9949 16355 10015 16356
rect 10501 16355 10567 16358
rect 12014 16356 12020 16358
rect 12084 16356 12090 16420
rect 8842 16352 9158 16353
rect 8842 16288 8848 16352
rect 8912 16288 8928 16352
rect 8992 16288 9008 16352
rect 9072 16288 9088 16352
rect 9152 16288 9158 16352
rect 8842 16287 9158 16288
rect 12790 16352 13106 16353
rect 12790 16288 12796 16352
rect 12860 16288 12876 16352
rect 12940 16288 12956 16352
rect 13020 16288 13036 16352
rect 13100 16288 13106 16352
rect 12790 16287 13106 16288
rect 7281 16280 7666 16282
rect 7281 16224 7286 16280
rect 7342 16224 7666 16280
rect 7281 16222 7666 16224
rect 8017 16282 8083 16285
rect 8477 16282 8543 16285
rect 8017 16280 8543 16282
rect 8017 16224 8022 16280
rect 8078 16224 8482 16280
rect 8538 16224 8543 16280
rect 8017 16222 8543 16224
rect 7281 16219 7347 16222
rect 8017 16219 8083 16222
rect 8477 16219 8543 16222
rect 9305 16282 9371 16285
rect 11697 16282 11763 16285
rect 9305 16280 11763 16282
rect 9305 16224 9310 16280
rect 9366 16224 11702 16280
rect 11758 16224 11763 16280
rect 9305 16222 11763 16224
rect 9305 16219 9371 16222
rect 11697 16219 11763 16222
rect 9765 16146 9831 16149
rect 13077 16146 13143 16149
rect 4340 16144 13143 16146
rect 4340 16088 9770 16144
rect 9826 16088 13082 16144
rect 13138 16088 13143 16144
rect 4340 16086 13143 16088
rect 9765 16083 9831 16086
rect 13077 16083 13143 16086
rect 2221 16010 2287 16013
rect 2446 16010 2452 16012
rect 2221 16008 2452 16010
rect 2221 15952 2226 16008
rect 2282 15952 2452 16008
rect 2221 15950 2452 15952
rect 2221 15947 2287 15950
rect 2446 15948 2452 15950
rect 2516 15948 2522 16012
rect 3969 16010 4035 16013
rect 11830 16010 11836 16012
rect 3969 16008 11836 16010
rect 3969 15952 3974 16008
rect 4030 15952 11836 16008
rect 3969 15950 11836 15952
rect 3969 15947 4035 15950
rect 11830 15948 11836 15950
rect 11900 15948 11906 16012
rect 4286 15812 4292 15876
rect 4356 15874 4362 15876
rect 5073 15874 5139 15877
rect 5390 15874 5396 15876
rect 4356 15872 5396 15874
rect 4356 15816 5078 15872
rect 5134 15816 5396 15872
rect 4356 15814 5396 15816
rect 4356 15812 4362 15814
rect 5073 15811 5139 15814
rect 5390 15812 5396 15814
rect 5460 15812 5466 15876
rect 7741 15874 7807 15877
rect 8702 15874 8708 15876
rect 7741 15872 8708 15874
rect 7741 15816 7746 15872
rect 7802 15816 8708 15872
rect 7741 15814 8708 15816
rect 7741 15811 7807 15814
rect 8702 15812 8708 15814
rect 8772 15874 8778 15876
rect 9029 15874 9095 15877
rect 8772 15872 9095 15874
rect 8772 15816 9034 15872
rect 9090 15816 9095 15872
rect 8772 15814 9095 15816
rect 8772 15812 8778 15814
rect 9029 15811 9095 15814
rect 9305 15874 9371 15877
rect 10593 15874 10659 15877
rect 9305 15872 10659 15874
rect 9305 15816 9310 15872
rect 9366 15816 10598 15872
rect 10654 15816 10659 15872
rect 9305 15814 10659 15816
rect 9305 15811 9371 15814
rect 10593 15811 10659 15814
rect 11513 15874 11579 15877
rect 13169 15874 13235 15877
rect 11513 15872 13235 15874
rect 11513 15816 11518 15872
rect 11574 15816 13174 15872
rect 13230 15816 13235 15872
rect 11513 15814 13235 15816
rect 11513 15811 11579 15814
rect 2920 15808 3236 15809
rect 0 15738 400 15768
rect 2920 15744 2926 15808
rect 2990 15744 3006 15808
rect 3070 15744 3086 15808
rect 3150 15744 3166 15808
rect 3230 15744 3236 15808
rect 2920 15743 3236 15744
rect 6868 15808 7184 15809
rect 6868 15744 6874 15808
rect 6938 15744 6954 15808
rect 7018 15744 7034 15808
rect 7098 15744 7114 15808
rect 7178 15744 7184 15808
rect 6868 15743 7184 15744
rect 10816 15808 11132 15809
rect 10816 15744 10822 15808
rect 10886 15744 10902 15808
rect 10966 15744 10982 15808
rect 11046 15744 11062 15808
rect 11126 15744 11132 15808
rect 10816 15743 11132 15744
rect 11700 15741 11760 15814
rect 13169 15811 13235 15814
rect 14764 15808 15080 15809
rect 14764 15744 14770 15808
rect 14834 15744 14850 15808
rect 14914 15744 14930 15808
rect 14994 15744 15010 15808
rect 15074 15744 15080 15808
rect 14764 15743 15080 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 400 15678
rect 1393 15675 1459 15678
rect 7276 15676 7282 15740
rect 7346 15738 7352 15740
rect 7966 15738 7972 15740
rect 7346 15678 7972 15738
rect 7346 15676 7352 15678
rect 7966 15676 7972 15678
rect 8036 15676 8042 15740
rect 10593 15738 10659 15741
rect 8158 15736 10659 15738
rect 8158 15680 10598 15736
rect 10654 15680 10659 15736
rect 8158 15678 10659 15680
rect 3550 15540 3556 15604
rect 3620 15602 3626 15604
rect 6269 15602 6335 15605
rect 8158 15602 8218 15678
rect 10593 15675 10659 15678
rect 11697 15736 11763 15741
rect 11697 15680 11702 15736
rect 11758 15680 11763 15736
rect 11697 15675 11763 15680
rect 12758 15678 14704 15738
rect 3620 15600 8218 15602
rect 3620 15544 6274 15600
rect 6330 15544 8218 15600
rect 3620 15542 8218 15544
rect 3620 15540 3626 15542
rect 6269 15539 6335 15542
rect 8334 15540 8340 15604
rect 8404 15602 8410 15604
rect 10777 15602 10843 15605
rect 8404 15600 10843 15602
rect 8404 15544 10782 15600
rect 10838 15544 10843 15600
rect 8404 15542 10843 15544
rect 8404 15540 8410 15542
rect 10777 15539 10843 15542
rect 10961 15602 11027 15605
rect 12758 15602 12818 15678
rect 10961 15600 12818 15602
rect 10961 15544 10966 15600
rect 11022 15544 12818 15600
rect 10961 15542 12818 15544
rect 12893 15602 12959 15605
rect 13721 15602 13787 15605
rect 12893 15600 13787 15602
rect 12893 15544 12898 15600
rect 12954 15544 13726 15600
rect 13782 15544 13787 15600
rect 12893 15542 13787 15544
rect 14644 15602 14704 15678
rect 15878 15602 15884 15604
rect 14644 15542 15884 15602
rect 10961 15539 11027 15542
rect 12893 15539 12959 15542
rect 13721 15539 13787 15542
rect 15878 15540 15884 15542
rect 15948 15540 15954 15604
rect 657 15466 723 15469
rect 8937 15466 9003 15469
rect 657 15464 9003 15466
rect 657 15408 662 15464
rect 718 15408 8942 15464
rect 8998 15408 9003 15464
rect 657 15406 9003 15408
rect 657 15403 723 15406
rect 8937 15403 9003 15406
rect 9213 15466 9279 15469
rect 9489 15466 9555 15469
rect 9213 15464 9555 15466
rect 9213 15408 9218 15464
rect 9274 15408 9494 15464
rect 9550 15408 9555 15464
rect 9213 15406 9555 15408
rect 9213 15403 9279 15406
rect 9489 15403 9555 15406
rect 9806 15404 9812 15468
rect 9876 15466 9882 15468
rect 12709 15466 12775 15469
rect 9876 15464 12775 15466
rect 9876 15408 12714 15464
rect 12770 15408 12775 15464
rect 9876 15406 12775 15408
rect 9876 15404 9882 15406
rect 12709 15403 12775 15406
rect 12985 15466 13051 15469
rect 13854 15466 13860 15468
rect 12985 15464 13860 15466
rect 12985 15408 12990 15464
rect 13046 15408 13860 15464
rect 12985 15406 13860 15408
rect 12985 15403 13051 15406
rect 13854 15404 13860 15406
rect 13924 15404 13930 15468
rect 1894 15268 1900 15332
rect 1964 15330 1970 15332
rect 4613 15330 4679 15333
rect 1964 15328 4679 15330
rect 1964 15272 4618 15328
rect 4674 15272 4679 15328
rect 1964 15270 4679 15272
rect 1964 15268 1970 15270
rect 4613 15267 4679 15270
rect 5390 15268 5396 15332
rect 5460 15330 5466 15332
rect 6637 15330 6703 15333
rect 5460 15328 6703 15330
rect 5460 15272 6642 15328
rect 6698 15272 6703 15328
rect 5460 15270 6703 15272
rect 5460 15268 5466 15270
rect 6637 15267 6703 15270
rect 7598 15268 7604 15332
rect 7668 15330 7674 15332
rect 10317 15330 10383 15333
rect 12157 15330 12223 15333
rect 7668 15270 8770 15330
rect 7668 15268 7674 15270
rect 4894 15264 5210 15265
rect 4894 15200 4900 15264
rect 4964 15200 4980 15264
rect 5044 15200 5060 15264
rect 5124 15200 5140 15264
rect 5204 15200 5210 15264
rect 4894 15199 5210 15200
rect 6085 15196 6151 15197
rect 6085 15194 6132 15196
rect 6040 15192 6132 15194
rect 6040 15136 6090 15192
rect 6040 15134 6132 15136
rect 6085 15132 6132 15134
rect 6196 15132 6202 15196
rect 6085 15131 6151 15132
rect 6126 14996 6132 15060
rect 6196 15058 6202 15060
rect 7189 15058 7255 15061
rect 7465 15058 7531 15061
rect 6196 15056 7531 15058
rect 6196 15000 7194 15056
rect 7250 15000 7470 15056
rect 7526 15000 7531 15056
rect 6196 14998 7531 15000
rect 8710 15058 8770 15270
rect 9262 15328 12223 15330
rect 9262 15272 10322 15328
rect 10378 15272 12162 15328
rect 12218 15272 12223 15328
rect 9262 15270 12223 15272
rect 8842 15264 9158 15265
rect 8842 15200 8848 15264
rect 8912 15200 8928 15264
rect 8992 15200 9008 15264
rect 9072 15200 9088 15264
rect 9152 15200 9158 15264
rect 8842 15199 9158 15200
rect 9262 15058 9322 15270
rect 10317 15267 10383 15270
rect 12157 15267 12223 15270
rect 12790 15264 13106 15265
rect 12790 15200 12796 15264
rect 12860 15200 12876 15264
rect 12940 15200 12956 15264
rect 13020 15200 13036 15264
rect 13100 15200 13106 15264
rect 12790 15199 13106 15200
rect 11053 15194 11119 15197
rect 11278 15194 11284 15196
rect 11053 15192 11284 15194
rect 11053 15136 11058 15192
rect 11114 15136 11284 15192
rect 11053 15134 11284 15136
rect 11053 15131 11119 15134
rect 11278 15132 11284 15134
rect 11348 15132 11354 15196
rect 12065 15194 12131 15197
rect 12382 15194 12388 15196
rect 12065 15192 12388 15194
rect 12065 15136 12070 15192
rect 12126 15136 12388 15192
rect 12065 15134 12388 15136
rect 12065 15131 12131 15134
rect 12382 15132 12388 15134
rect 12452 15132 12458 15196
rect 8710 14998 9322 15058
rect 6196 14996 6202 14998
rect 7189 14995 7255 14998
rect 7465 14995 7531 14998
rect 9806 14996 9812 15060
rect 9876 15058 9882 15060
rect 9949 15058 10015 15061
rect 9876 15056 10015 15058
rect 9876 15000 9954 15056
rect 10010 15000 10015 15056
rect 9876 14998 10015 15000
rect 9876 14996 9882 14998
rect 9949 14995 10015 14998
rect 10174 14996 10180 15060
rect 10244 15058 10250 15060
rect 10501 15058 10567 15061
rect 10244 15056 10567 15058
rect 10244 15000 10506 15056
rect 10562 15000 10567 15056
rect 10244 14998 10567 15000
rect 10244 14996 10250 14998
rect 10501 14995 10567 14998
rect 11605 15058 11671 15061
rect 15510 15058 15516 15060
rect 11605 15056 15516 15058
rect 11605 15000 11610 15056
rect 11666 15000 15516 15056
rect 11605 14998 15516 15000
rect 11605 14995 11671 14998
rect 15510 14996 15516 14998
rect 15580 14996 15586 15060
rect 3734 14922 3740 14924
rect 3558 14862 3740 14922
rect 2920 14720 3236 14721
rect 2920 14656 2926 14720
rect 2990 14656 3006 14720
rect 3070 14656 3086 14720
rect 3150 14656 3166 14720
rect 3230 14656 3236 14720
rect 2920 14655 3236 14656
rect 2262 14588 2268 14652
rect 2332 14650 2338 14652
rect 2589 14650 2655 14653
rect 2332 14648 2655 14650
rect 2332 14592 2594 14648
rect 2650 14592 2655 14648
rect 2332 14590 2655 14592
rect 3558 14650 3618 14862
rect 3734 14860 3740 14862
rect 3804 14860 3810 14924
rect 4470 14860 4476 14924
rect 4540 14922 4546 14924
rect 4889 14922 4955 14925
rect 4540 14920 4955 14922
rect 4540 14864 4894 14920
rect 4950 14864 4955 14920
rect 4540 14862 4955 14864
rect 4540 14860 4546 14862
rect 4889 14859 4955 14862
rect 6453 14922 6519 14925
rect 8477 14922 8543 14925
rect 9305 14922 9371 14925
rect 12065 14922 12131 14925
rect 6453 14920 7896 14922
rect 6453 14864 6458 14920
rect 6514 14864 7896 14920
rect 6453 14862 7896 14864
rect 6453 14859 6519 14862
rect 3734 14724 3740 14788
rect 3804 14786 3810 14788
rect 6456 14786 6516 14859
rect 3804 14726 6516 14786
rect 3804 14724 3810 14726
rect 6868 14720 7184 14721
rect 6868 14656 6874 14720
rect 6938 14656 6954 14720
rect 7018 14656 7034 14720
rect 7098 14656 7114 14720
rect 7178 14656 7184 14720
rect 6868 14655 7184 14656
rect 4521 14652 4587 14653
rect 4470 14650 4476 14652
rect 3558 14590 3802 14650
rect 4430 14590 4476 14650
rect 4540 14648 4587 14652
rect 4582 14592 4587 14648
rect 2332 14588 2338 14590
rect 2589 14587 2655 14590
rect 2262 14316 2268 14380
rect 2332 14378 2338 14380
rect 3550 14378 3556 14380
rect 2332 14318 3556 14378
rect 2332 14316 2338 14318
rect 3550 14316 3556 14318
rect 3620 14316 3626 14380
rect 0 14242 400 14272
rect 1485 14242 1551 14245
rect 0 14240 1551 14242
rect 0 14184 1490 14240
rect 1546 14184 1551 14240
rect 0 14182 1551 14184
rect 0 14152 400 14182
rect 1485 14179 1551 14182
rect 3550 14180 3556 14244
rect 3620 14242 3626 14244
rect 3742 14242 3802 14590
rect 4470 14588 4476 14590
rect 4540 14588 4587 14592
rect 4521 14587 4587 14588
rect 6177 14650 6243 14653
rect 6729 14650 6795 14653
rect 6177 14648 6795 14650
rect 6177 14592 6182 14648
rect 6238 14592 6734 14648
rect 6790 14592 6795 14648
rect 6177 14590 6795 14592
rect 7836 14650 7896 14862
rect 8477 14920 9371 14922
rect 8477 14864 8482 14920
rect 8538 14864 9310 14920
rect 9366 14864 9371 14920
rect 8477 14862 9371 14864
rect 8477 14859 8543 14862
rect 9305 14859 9371 14862
rect 10596 14920 12131 14922
rect 10596 14864 12070 14920
rect 12126 14864 12131 14920
rect 10596 14862 12131 14864
rect 7966 14724 7972 14788
rect 8036 14786 8042 14788
rect 9121 14786 9187 14789
rect 8036 14784 9187 14786
rect 8036 14728 9126 14784
rect 9182 14728 9187 14784
rect 8036 14726 9187 14728
rect 8036 14724 8042 14726
rect 9121 14723 9187 14726
rect 9254 14724 9260 14788
rect 9324 14786 9330 14788
rect 10596 14786 10656 14862
rect 12065 14859 12131 14862
rect 12617 14922 12683 14925
rect 16430 14922 16436 14924
rect 12617 14920 16436 14922
rect 12617 14864 12622 14920
rect 12678 14864 16436 14920
rect 12617 14862 16436 14864
rect 12617 14859 12683 14862
rect 16430 14860 16436 14862
rect 16500 14860 16506 14924
rect 9324 14726 10656 14786
rect 13537 14786 13603 14789
rect 13670 14786 13676 14788
rect 13537 14784 13676 14786
rect 13537 14728 13542 14784
rect 13598 14728 13676 14784
rect 13537 14726 13676 14728
rect 9324 14724 9330 14726
rect 13537 14723 13603 14726
rect 13670 14724 13676 14726
rect 13740 14724 13746 14788
rect 10816 14720 11132 14721
rect 10816 14656 10822 14720
rect 10886 14656 10902 14720
rect 10966 14656 10982 14720
rect 11046 14656 11062 14720
rect 11126 14656 11132 14720
rect 10816 14655 11132 14656
rect 14764 14720 15080 14721
rect 14764 14656 14770 14720
rect 14834 14656 14850 14720
rect 14914 14656 14930 14720
rect 14994 14656 15010 14720
rect 15074 14656 15080 14720
rect 14764 14655 15080 14656
rect 10501 14650 10567 14653
rect 7836 14648 10567 14650
rect 7836 14592 10506 14648
rect 10562 14592 10567 14648
rect 7836 14590 10567 14592
rect 6177 14587 6243 14590
rect 6729 14587 6795 14590
rect 10501 14587 10567 14590
rect 12198 14588 12204 14652
rect 12268 14650 12274 14652
rect 12709 14650 12775 14653
rect 12268 14648 12775 14650
rect 12268 14592 12714 14648
rect 12770 14592 12775 14648
rect 12268 14590 12775 14592
rect 12268 14588 12274 14590
rect 12709 14587 12775 14590
rect 4797 14514 4863 14517
rect 5349 14514 5415 14517
rect 4797 14512 5415 14514
rect 4797 14456 4802 14512
rect 4858 14456 5354 14512
rect 5410 14456 5415 14512
rect 4797 14454 5415 14456
rect 4797 14451 4863 14454
rect 5349 14451 5415 14454
rect 6453 14514 6519 14517
rect 7465 14514 7531 14517
rect 8753 14514 8819 14517
rect 6453 14512 7531 14514
rect 6453 14456 6458 14512
rect 6514 14456 7470 14512
rect 7526 14456 7531 14512
rect 6453 14454 7531 14456
rect 6453 14451 6519 14454
rect 7465 14451 7531 14454
rect 8250 14512 8819 14514
rect 8250 14456 8758 14512
rect 8814 14456 8819 14512
rect 8250 14454 8819 14456
rect 3918 14316 3924 14380
rect 3988 14378 3994 14380
rect 4429 14378 4495 14381
rect 8250 14378 8310 14454
rect 8753 14451 8819 14454
rect 9121 14514 9187 14517
rect 10777 14514 10843 14517
rect 9121 14512 10843 14514
rect 9121 14456 9126 14512
rect 9182 14456 10782 14512
rect 10838 14456 10843 14512
rect 9121 14454 10843 14456
rect 9121 14451 9187 14454
rect 10777 14451 10843 14454
rect 10961 14514 11027 14517
rect 11881 14514 11947 14517
rect 13537 14516 13603 14517
rect 13486 14514 13492 14516
rect 10961 14512 11947 14514
rect 10961 14456 10966 14512
rect 11022 14456 11886 14512
rect 11942 14456 11947 14512
rect 10961 14454 11947 14456
rect 13446 14454 13492 14514
rect 13556 14512 13603 14516
rect 13598 14456 13603 14512
rect 10961 14451 11027 14454
rect 11881 14451 11947 14454
rect 13486 14452 13492 14454
rect 13556 14452 13603 14456
rect 13537 14451 13603 14452
rect 3988 14376 8310 14378
rect 3988 14320 4434 14376
rect 4490 14320 8310 14376
rect 3988 14318 8310 14320
rect 8710 14318 9322 14378
rect 3988 14316 3994 14318
rect 4429 14315 4495 14318
rect 3620 14182 3802 14242
rect 4061 14240 4127 14245
rect 4061 14184 4066 14240
rect 4122 14184 4127 14240
rect 3620 14180 3626 14182
rect 4061 14179 4127 14184
rect 6729 14242 6795 14245
rect 8569 14242 8635 14245
rect 6729 14240 8635 14242
rect 6729 14184 6734 14240
rect 6790 14184 8574 14240
rect 8630 14184 8635 14240
rect 6729 14182 8635 14184
rect 6729 14179 6795 14182
rect 8569 14179 8635 14182
rect 4064 14106 4124 14179
rect 4894 14176 5210 14177
rect 4894 14112 4900 14176
rect 4964 14112 4980 14176
rect 5044 14112 5060 14176
rect 5124 14112 5140 14176
rect 5204 14112 5210 14176
rect 4894 14111 5210 14112
rect 3328 14046 4124 14106
rect 749 13834 815 13837
rect 2957 13834 3023 13837
rect 749 13832 3023 13834
rect 749 13776 754 13832
rect 810 13776 2962 13832
rect 3018 13776 3023 13832
rect 749 13774 3023 13776
rect 749 13771 815 13774
rect 2957 13771 3023 13774
rect 2920 13632 3236 13633
rect 2920 13568 2926 13632
rect 2990 13568 3006 13632
rect 3070 13568 3086 13632
rect 3150 13568 3166 13632
rect 3230 13568 3236 13632
rect 2920 13567 3236 13568
rect 1577 13426 1643 13429
rect 1853 13426 1919 13429
rect 2865 13426 2931 13429
rect 1577 13424 2931 13426
rect 1577 13368 1582 13424
rect 1638 13368 1858 13424
rect 1914 13368 2870 13424
rect 2926 13368 2931 13424
rect 1577 13366 2931 13368
rect 1577 13363 1643 13366
rect 1853 13363 1919 13366
rect 2865 13363 2931 13366
rect 3141 13426 3207 13429
rect 3328 13426 3388 14046
rect 5942 14044 5948 14108
rect 6012 14106 6018 14108
rect 8710 14106 8770 14318
rect 8842 14176 9158 14177
rect 8842 14112 8848 14176
rect 8912 14112 8928 14176
rect 8992 14112 9008 14176
rect 9072 14112 9088 14176
rect 9152 14112 9158 14176
rect 8842 14111 9158 14112
rect 6012 14046 8770 14106
rect 9262 14106 9322 14318
rect 9622 14316 9628 14380
rect 9692 14378 9698 14380
rect 14917 14378 14983 14381
rect 9692 14376 14983 14378
rect 9692 14320 14922 14376
rect 14978 14320 14983 14376
rect 9692 14318 14983 14320
rect 9692 14316 9698 14318
rect 14917 14315 14983 14318
rect 9397 14242 9463 14245
rect 10358 14242 10364 14244
rect 9397 14240 10364 14242
rect 9397 14184 9402 14240
rect 9458 14184 10364 14240
rect 9397 14182 10364 14184
rect 9397 14179 9463 14182
rect 10358 14180 10364 14182
rect 10428 14180 10434 14244
rect 11278 14180 11284 14244
rect 11348 14242 11354 14244
rect 12157 14242 12223 14245
rect 11348 14240 12223 14242
rect 11348 14184 12162 14240
rect 12218 14184 12223 14240
rect 11348 14182 12223 14184
rect 11348 14180 11354 14182
rect 12157 14179 12223 14182
rect 13302 14180 13308 14244
rect 13372 14242 13378 14244
rect 13445 14242 13511 14245
rect 13372 14240 13511 14242
rect 13372 14184 13450 14240
rect 13506 14184 13511 14240
rect 13372 14182 13511 14184
rect 13372 14180 13378 14182
rect 13445 14179 13511 14182
rect 12790 14176 13106 14177
rect 12790 14112 12796 14176
rect 12860 14112 12876 14176
rect 12940 14112 12956 14176
rect 13020 14112 13036 14176
rect 13100 14112 13106 14176
rect 12790 14111 13106 14112
rect 11605 14106 11671 14109
rect 9262 14104 11671 14106
rect 9262 14048 11610 14104
rect 11666 14048 11671 14104
rect 9262 14046 11671 14048
rect 6012 14044 6018 14046
rect 11605 14043 11671 14046
rect 11789 14106 11855 14109
rect 12065 14106 12131 14109
rect 13997 14106 14063 14109
rect 11789 14104 12131 14106
rect 11789 14048 11794 14104
rect 11850 14048 12070 14104
rect 12126 14048 12131 14104
rect 11789 14046 12131 14048
rect 11789 14043 11855 14046
rect 12065 14043 12131 14046
rect 13494 14104 14063 14106
rect 13494 14048 14002 14104
rect 14058 14048 14063 14104
rect 13494 14046 14063 14048
rect 3969 13970 4035 13973
rect 13494 13970 13554 14046
rect 13997 14043 14063 14046
rect 3969 13968 13554 13970
rect 3969 13912 3974 13968
rect 4030 13912 13554 13968
rect 3969 13910 13554 13912
rect 13997 13970 14063 13973
rect 14406 13970 14412 13972
rect 13997 13968 14412 13970
rect 13997 13912 14002 13968
rect 14058 13912 14412 13968
rect 13997 13910 14412 13912
rect 3969 13907 4035 13910
rect 13997 13907 14063 13910
rect 14406 13908 14412 13910
rect 14476 13908 14482 13972
rect 4889 13834 4955 13837
rect 7741 13834 7807 13837
rect 4889 13832 7807 13834
rect 4889 13776 4894 13832
rect 4950 13776 7746 13832
rect 7802 13776 7807 13832
rect 4889 13774 7807 13776
rect 4889 13771 4955 13774
rect 7741 13771 7807 13774
rect 8702 13772 8708 13836
rect 8772 13834 8778 13836
rect 8845 13834 8911 13837
rect 12709 13834 12775 13837
rect 13445 13834 13511 13837
rect 8772 13832 13511 13834
rect 8772 13776 8850 13832
rect 8906 13776 12714 13832
rect 12770 13776 13450 13832
rect 13506 13776 13511 13832
rect 8772 13774 13511 13776
rect 8772 13772 8778 13774
rect 8845 13771 8911 13774
rect 12709 13771 12775 13774
rect 13445 13771 13511 13774
rect 13905 13834 13971 13837
rect 14549 13834 14615 13837
rect 13905 13832 14615 13834
rect 13905 13776 13910 13832
rect 13966 13776 14554 13832
rect 14610 13776 14615 13832
rect 13905 13774 14615 13776
rect 13905 13771 13971 13774
rect 14549 13771 14615 13774
rect 15101 13834 15167 13837
rect 15101 13832 15348 13834
rect 15101 13776 15106 13832
rect 15162 13776 15348 13832
rect 15101 13774 15348 13776
rect 15101 13771 15167 13774
rect 15288 13701 15348 13774
rect 4470 13636 4476 13700
rect 4540 13698 4546 13700
rect 4705 13698 4771 13701
rect 5625 13700 5691 13701
rect 5574 13698 5580 13700
rect 4540 13696 4771 13698
rect 4540 13640 4710 13696
rect 4766 13640 4771 13696
rect 4540 13638 4771 13640
rect 5534 13638 5580 13698
rect 5644 13696 5691 13700
rect 8937 13698 9003 13701
rect 9857 13698 9923 13701
rect 5686 13640 5691 13696
rect 4540 13636 4546 13638
rect 4705 13635 4771 13638
rect 5574 13636 5580 13638
rect 5644 13636 5691 13640
rect 5625 13635 5691 13636
rect 7284 13638 8632 13698
rect 6868 13632 7184 13633
rect 6868 13568 6874 13632
rect 6938 13568 6954 13632
rect 7018 13568 7034 13632
rect 7098 13568 7114 13632
rect 7178 13568 7184 13632
rect 6868 13567 7184 13568
rect 3877 13562 3943 13565
rect 5574 13562 5580 13564
rect 3877 13560 5580 13562
rect 3877 13504 3882 13560
rect 3938 13504 5580 13560
rect 3877 13502 5580 13504
rect 3877 13499 3943 13502
rect 5574 13500 5580 13502
rect 5644 13500 5650 13564
rect 7284 13528 7344 13638
rect 7238 13468 7344 13528
rect 7782 13500 7788 13564
rect 7852 13562 7858 13564
rect 8201 13562 8267 13565
rect 7852 13560 8267 13562
rect 7852 13504 8206 13560
rect 8262 13504 8267 13560
rect 7852 13502 8267 13504
rect 7852 13500 7858 13502
rect 8201 13499 8267 13502
rect 4521 13428 4587 13429
rect 3141 13424 3388 13426
rect 3141 13368 3146 13424
rect 3202 13368 3388 13424
rect 3141 13366 3388 13368
rect 3141 13363 3207 13366
rect 4470 13364 4476 13428
rect 4540 13426 4587 13428
rect 5809 13426 5875 13429
rect 7238 13426 7298 13468
rect 4540 13424 4632 13426
rect 4582 13368 4632 13424
rect 4540 13366 4632 13368
rect 5809 13424 7298 13426
rect 5809 13368 5814 13424
rect 5870 13368 7298 13424
rect 5809 13366 7298 13368
rect 8572 13426 8632 13638
rect 8937 13696 9923 13698
rect 8937 13640 8942 13696
rect 8998 13640 9862 13696
rect 9918 13640 9923 13696
rect 8937 13638 9923 13640
rect 8937 13635 9003 13638
rect 9857 13635 9923 13638
rect 11278 13636 11284 13700
rect 11348 13698 11354 13700
rect 12065 13698 12131 13701
rect 11348 13696 12131 13698
rect 11348 13640 12070 13696
rect 12126 13640 12131 13696
rect 11348 13638 12131 13640
rect 11348 13636 11354 13638
rect 12065 13635 12131 13638
rect 13997 13698 14063 13701
rect 14181 13698 14247 13701
rect 13997 13696 14247 13698
rect 13997 13640 14002 13696
rect 14058 13640 14186 13696
rect 14242 13640 14247 13696
rect 13997 13638 14247 13640
rect 13997 13635 14063 13638
rect 14181 13635 14247 13638
rect 14457 13698 14523 13701
rect 14590 13698 14596 13700
rect 14457 13696 14596 13698
rect 14457 13640 14462 13696
rect 14518 13640 14596 13696
rect 14457 13638 14596 13640
rect 14457 13635 14523 13638
rect 14590 13636 14596 13638
rect 14660 13636 14666 13700
rect 15285 13696 15351 13701
rect 15285 13640 15290 13696
rect 15346 13640 15351 13696
rect 15285 13635 15351 13640
rect 10816 13632 11132 13633
rect 10816 13568 10822 13632
rect 10886 13568 10902 13632
rect 10966 13568 10982 13632
rect 11046 13568 11062 13632
rect 11126 13568 11132 13632
rect 10816 13567 11132 13568
rect 14764 13632 15080 13633
rect 14764 13568 14770 13632
rect 14834 13568 14850 13632
rect 14914 13568 14930 13632
rect 14994 13568 15010 13632
rect 15074 13568 15080 13632
rect 14764 13567 15080 13568
rect 8702 13500 8708 13564
rect 8772 13562 8778 13564
rect 9121 13562 9187 13565
rect 8772 13560 9187 13562
rect 8772 13504 9126 13560
rect 9182 13504 9187 13560
rect 8772 13502 9187 13504
rect 8772 13500 8778 13502
rect 9121 13499 9187 13502
rect 11329 13562 11395 13565
rect 12985 13562 13051 13565
rect 11329 13560 13051 13562
rect 11329 13504 11334 13560
rect 11390 13504 12990 13560
rect 13046 13504 13051 13560
rect 11329 13502 13051 13504
rect 11329 13499 11395 13502
rect 12985 13499 13051 13502
rect 13164 13500 13170 13564
rect 13234 13562 13240 13564
rect 13537 13562 13603 13565
rect 13234 13560 13603 13562
rect 13234 13504 13542 13560
rect 13598 13504 13603 13560
rect 13234 13502 13603 13504
rect 13234 13500 13240 13502
rect 13537 13499 13603 13502
rect 13721 13562 13787 13565
rect 15377 13564 15443 13565
rect 14222 13562 14228 13564
rect 13721 13560 14228 13562
rect 13721 13504 13726 13560
rect 13782 13504 14228 13560
rect 13721 13502 14228 13504
rect 13721 13499 13787 13502
rect 14222 13500 14228 13502
rect 14292 13500 14298 13564
rect 15326 13500 15332 13564
rect 15396 13562 15443 13564
rect 15396 13560 15488 13562
rect 15438 13504 15488 13560
rect 15396 13502 15488 13504
rect 15396 13500 15443 13502
rect 15377 13499 15443 13500
rect 15377 13426 15443 13429
rect 8572 13424 15443 13426
rect 8572 13368 15382 13424
rect 15438 13368 15443 13424
rect 8572 13366 15443 13368
rect 4540 13364 4587 13366
rect 4521 13363 4587 13364
rect 5809 13363 5875 13366
rect 15377 13363 15443 13366
rect 2405 13290 2471 13293
rect 4521 13290 4587 13293
rect 4889 13290 4955 13293
rect 2405 13288 4955 13290
rect 2405 13232 2410 13288
rect 2466 13232 4526 13288
rect 4582 13232 4894 13288
rect 4950 13232 4955 13288
rect 2405 13230 4955 13232
rect 2405 13227 2471 13230
rect 4521 13227 4587 13230
rect 4889 13227 4955 13230
rect 6361 13290 6427 13293
rect 12157 13290 12223 13293
rect 6361 13288 12223 13290
rect 6361 13232 6366 13288
rect 6422 13232 12162 13288
rect 12218 13232 12223 13288
rect 6361 13230 12223 13232
rect 6361 13227 6427 13230
rect 12157 13227 12223 13230
rect 12525 13290 12591 13293
rect 15653 13292 15719 13293
rect 15142 13290 15148 13292
rect 12525 13288 15148 13290
rect 12525 13232 12530 13288
rect 12586 13232 15148 13288
rect 12525 13230 15148 13232
rect 12525 13227 12634 13230
rect 15142 13228 15148 13230
rect 15212 13228 15218 13292
rect 15653 13288 15700 13292
rect 15764 13290 15770 13292
rect 15653 13232 15658 13288
rect 15653 13228 15700 13232
rect 15764 13230 15810 13290
rect 15764 13228 15770 13230
rect 15653 13227 15719 13228
rect 3877 13154 3943 13157
rect 4061 13154 4127 13157
rect 3877 13152 4127 13154
rect 3877 13096 3882 13152
rect 3938 13096 4066 13152
rect 4122 13096 4127 13152
rect 3877 13094 4127 13096
rect 3877 13091 3943 13094
rect 4061 13091 4127 13094
rect 5809 13154 5875 13157
rect 5942 13154 5948 13156
rect 5809 13152 5948 13154
rect 5809 13096 5814 13152
rect 5870 13096 5948 13152
rect 5809 13094 5948 13096
rect 5809 13091 5875 13094
rect 5942 13092 5948 13094
rect 6012 13092 6018 13156
rect 6637 13154 6703 13157
rect 9489 13154 9555 13157
rect 11421 13154 11487 13157
rect 6637 13152 7068 13154
rect 6637 13096 6642 13152
rect 6698 13096 7068 13152
rect 6637 13094 7068 13096
rect 6637 13091 6703 13094
rect 4894 13088 5210 13089
rect 4894 13024 4900 13088
rect 4964 13024 4980 13088
rect 5044 13024 5060 13088
rect 5124 13024 5140 13088
rect 5204 13024 5210 13088
rect 4894 13023 5210 13024
rect 7008 13021 7068 13094
rect 9489 13152 11487 13154
rect 9489 13096 9494 13152
rect 9550 13096 11426 13152
rect 11482 13096 11487 13152
rect 9489 13094 11487 13096
rect 9489 13091 9555 13094
rect 11421 13091 11487 13094
rect 11646 13092 11652 13156
rect 11716 13154 11722 13156
rect 12433 13154 12499 13157
rect 11716 13152 12499 13154
rect 11716 13096 12438 13152
rect 12494 13096 12499 13152
rect 11716 13094 12499 13096
rect 11716 13092 11722 13094
rect 12433 13091 12499 13094
rect 8842 13088 9158 13089
rect 8842 13024 8848 13088
rect 8912 13024 8928 13088
rect 8992 13024 9008 13088
rect 9072 13024 9088 13088
rect 9152 13024 9158 13088
rect 8842 13023 9158 13024
rect 1577 13018 1643 13021
rect 4705 13020 4771 13021
rect 3734 13018 3740 13020
rect 1577 13016 3740 13018
rect 1577 12960 1582 13016
rect 1638 12960 3740 13016
rect 1577 12958 3740 12960
rect 1577 12955 1643 12958
rect 3734 12956 3740 12958
rect 3804 12956 3810 13020
rect 4654 12956 4660 13020
rect 4724 13018 4771 13020
rect 6177 13018 6243 13021
rect 4724 13016 4816 13018
rect 4766 12960 4816 13016
rect 4724 12958 4816 12960
rect 6177 13016 6562 13018
rect 6177 12960 6182 13016
rect 6238 12960 6562 13016
rect 6177 12958 6562 12960
rect 4724 12956 4771 12958
rect 4705 12955 4771 12956
rect 6177 12955 6243 12958
rect 2221 12880 2287 12885
rect 2221 12824 2226 12880
rect 2282 12824 2287 12880
rect 2221 12819 2287 12824
rect 3550 12820 3556 12884
rect 3620 12882 3626 12884
rect 3918 12882 3924 12884
rect 3620 12822 3924 12882
rect 3620 12820 3626 12822
rect 3918 12820 3924 12822
rect 3988 12820 3994 12884
rect 6126 12820 6132 12884
rect 6196 12882 6202 12884
rect 6361 12882 6427 12885
rect 6196 12880 6427 12882
rect 6196 12824 6366 12880
rect 6422 12824 6427 12880
rect 6196 12822 6427 12824
rect 6196 12820 6202 12822
rect 6361 12819 6427 12822
rect 0 12746 400 12776
rect 1945 12746 2011 12749
rect 0 12744 2011 12746
rect 0 12688 1950 12744
rect 2006 12688 2011 12744
rect 0 12686 2011 12688
rect 2224 12746 2284 12819
rect 3693 12746 3759 12749
rect 2224 12744 3759 12746
rect 2224 12688 3698 12744
rect 3754 12688 3759 12744
rect 2224 12686 3759 12688
rect 0 12656 400 12686
rect 1945 12683 2011 12686
rect 3693 12683 3759 12686
rect 4654 12684 4660 12748
rect 4724 12746 4730 12748
rect 4889 12746 4955 12749
rect 4724 12744 4955 12746
rect 4724 12688 4894 12744
rect 4950 12688 4955 12744
rect 4724 12686 4955 12688
rect 4724 12684 4730 12686
rect 4889 12683 4955 12686
rect 5441 12746 5507 12749
rect 5758 12746 5764 12748
rect 5441 12744 5764 12746
rect 5441 12688 5446 12744
rect 5502 12688 5764 12744
rect 5441 12686 5764 12688
rect 5441 12683 5507 12686
rect 5758 12684 5764 12686
rect 5828 12684 5834 12748
rect 6361 12746 6427 12749
rect 6502 12746 6562 12958
rect 7005 13016 7071 13021
rect 7005 12960 7010 13016
rect 7066 12960 7071 13016
rect 7005 12955 7071 12960
rect 7741 13018 7807 13021
rect 8150 13018 8156 13020
rect 7741 13016 8156 13018
rect 7741 12960 7746 13016
rect 7802 12960 8156 13016
rect 7741 12958 8156 12960
rect 7741 12955 7807 12958
rect 8150 12956 8156 12958
rect 8220 12956 8226 13020
rect 8477 13018 8543 13021
rect 8661 13018 8727 13021
rect 8477 13016 8727 13018
rect 8477 12960 8482 13016
rect 8538 12960 8666 13016
rect 8722 12960 8727 13016
rect 8477 12958 8727 12960
rect 8477 12955 8543 12958
rect 8661 12955 8727 12958
rect 9949 13018 10015 13021
rect 11329 13018 11395 13021
rect 9949 13016 11395 13018
rect 9949 12960 9954 13016
rect 10010 12960 11334 13016
rect 11390 12960 11395 13016
rect 9949 12958 11395 12960
rect 9949 12955 10015 12958
rect 11329 12955 11395 12958
rect 11513 13018 11579 13021
rect 11646 13018 11652 13020
rect 11513 13016 11652 13018
rect 11513 12960 11518 13016
rect 11574 12960 11652 13016
rect 11513 12958 11652 12960
rect 11513 12955 11579 12958
rect 11646 12956 11652 12958
rect 11716 12956 11722 13020
rect 12433 13018 12499 13021
rect 12574 13018 12634 13227
rect 17493 13154 17559 13157
rect 13172 13152 17559 13154
rect 13172 13096 17498 13152
rect 17554 13096 17559 13152
rect 13172 13094 17559 13096
rect 12790 13088 13106 13089
rect 12790 13024 12796 13088
rect 12860 13024 12876 13088
rect 12940 13024 12956 13088
rect 13020 13024 13036 13088
rect 13100 13024 13106 13088
rect 12790 13023 13106 13024
rect 12433 13016 12634 13018
rect 12433 12960 12438 13016
rect 12494 12960 12634 13016
rect 12433 12958 12634 12960
rect 12433 12955 12499 12958
rect 7373 12882 7439 12885
rect 6870 12880 7439 12882
rect 6870 12824 7378 12880
rect 7434 12824 7439 12880
rect 6870 12822 7439 12824
rect 6870 12746 6930 12822
rect 7373 12819 7439 12822
rect 7557 12882 7623 12885
rect 13172 12882 13232 13094
rect 17493 13091 17559 13094
rect 13445 13018 13511 13021
rect 14181 13018 14247 13021
rect 13445 13016 14247 13018
rect 13445 12960 13450 13016
rect 13506 12960 14186 13016
rect 14242 12960 14247 13016
rect 13445 12958 14247 12960
rect 13445 12955 13511 12958
rect 14181 12955 14247 12958
rect 14365 13018 14431 13021
rect 16062 13018 16068 13020
rect 14365 13016 16068 13018
rect 14365 12960 14370 13016
rect 14426 12960 16068 13016
rect 14365 12958 16068 12960
rect 14365 12955 14431 12958
rect 16062 12956 16068 12958
rect 16132 12956 16138 13020
rect 13813 12882 13879 12885
rect 7557 12880 12634 12882
rect 7557 12824 7562 12880
rect 7618 12848 12634 12880
rect 12712 12848 13232 12882
rect 7618 12824 13232 12848
rect 7557 12822 13232 12824
rect 13310 12880 13879 12882
rect 13310 12824 13818 12880
rect 13874 12824 13879 12880
rect 13310 12822 13879 12824
rect 7557 12819 7623 12822
rect 12574 12788 12772 12822
rect 6361 12744 6562 12746
rect 6361 12688 6366 12744
rect 6422 12688 6562 12744
rect 6361 12686 6562 12688
rect 6732 12686 6930 12746
rect 7005 12746 7071 12749
rect 7741 12746 7807 12749
rect 7005 12744 7807 12746
rect 7005 12688 7010 12744
rect 7066 12688 7746 12744
rect 7802 12688 7807 12744
rect 7005 12686 7807 12688
rect 6361 12683 6427 12686
rect 3601 12612 3667 12613
rect 3550 12610 3556 12612
rect 3510 12550 3556 12610
rect 3620 12608 3667 12612
rect 3662 12552 3667 12608
rect 3550 12548 3556 12550
rect 3620 12548 3667 12552
rect 3734 12548 3740 12612
rect 3804 12610 3810 12612
rect 4337 12610 4403 12613
rect 3804 12608 4403 12610
rect 3804 12552 4342 12608
rect 4398 12552 4403 12608
rect 3804 12550 4403 12552
rect 3804 12548 3810 12550
rect 3601 12547 3667 12548
rect 4337 12547 4403 12550
rect 5165 12610 5231 12613
rect 6732 12610 6792 12686
rect 7005 12683 7071 12686
rect 7741 12683 7807 12686
rect 7925 12746 7991 12749
rect 9121 12746 9187 12749
rect 7925 12744 9187 12746
rect 7925 12688 7930 12744
rect 7986 12688 9126 12744
rect 9182 12688 9187 12744
rect 7925 12686 9187 12688
rect 7925 12683 7991 12686
rect 9121 12683 9187 12686
rect 9438 12684 9444 12748
rect 9508 12746 9514 12748
rect 9765 12746 9831 12749
rect 12433 12746 12499 12749
rect 9508 12744 9831 12746
rect 9508 12688 9770 12744
rect 9826 12688 9831 12744
rect 9508 12686 9831 12688
rect 9508 12684 9514 12686
rect 9765 12683 9831 12686
rect 10688 12744 12499 12746
rect 10688 12688 12438 12744
rect 12494 12688 12499 12744
rect 10688 12686 12499 12688
rect 5165 12608 6792 12610
rect 5165 12552 5170 12608
rect 5226 12552 6792 12608
rect 5165 12550 6792 12552
rect 7465 12610 7531 12613
rect 7782 12610 7788 12612
rect 7465 12608 7788 12610
rect 7465 12552 7470 12608
rect 7526 12552 7788 12608
rect 7465 12550 7788 12552
rect 5165 12547 5231 12550
rect 7465 12547 7531 12550
rect 7782 12548 7788 12550
rect 7852 12548 7858 12612
rect 8017 12610 8083 12613
rect 8150 12610 8156 12612
rect 8017 12608 8156 12610
rect 8017 12552 8022 12608
rect 8078 12552 8156 12608
rect 8017 12550 8156 12552
rect 8017 12547 8083 12550
rect 8150 12548 8156 12550
rect 8220 12548 8226 12612
rect 9438 12548 9444 12612
rect 9508 12610 9514 12612
rect 10225 12610 10291 12613
rect 9508 12608 10291 12610
rect 9508 12552 10230 12608
rect 10286 12552 10291 12608
rect 9508 12550 10291 12552
rect 9508 12548 9514 12550
rect 10225 12547 10291 12550
rect 2920 12544 3236 12545
rect 2920 12480 2926 12544
rect 2990 12480 3006 12544
rect 3070 12480 3086 12544
rect 3150 12480 3166 12544
rect 3230 12480 3236 12544
rect 2920 12479 3236 12480
rect 6868 12544 7184 12545
rect 6868 12480 6874 12544
rect 6938 12480 6954 12544
rect 7018 12480 7034 12544
rect 7098 12480 7114 12544
rect 7178 12480 7184 12544
rect 6868 12479 7184 12480
rect 4286 12412 4292 12476
rect 4356 12474 4362 12476
rect 4521 12474 4587 12477
rect 4356 12472 4587 12474
rect 4356 12416 4526 12472
rect 4582 12416 4587 12472
rect 4356 12414 4587 12416
rect 4356 12412 4362 12414
rect 4521 12411 4587 12414
rect 4797 12474 4863 12477
rect 6494 12474 6500 12476
rect 4797 12472 6500 12474
rect 4797 12416 4802 12472
rect 4858 12416 6500 12472
rect 4797 12414 6500 12416
rect 4797 12411 4863 12414
rect 6494 12412 6500 12414
rect 6564 12412 6570 12476
rect 8702 12474 8708 12476
rect 7744 12414 8708 12474
rect 2589 12338 2655 12341
rect 4286 12338 4292 12340
rect 2589 12336 4292 12338
rect 2589 12280 2594 12336
rect 2650 12280 4292 12336
rect 2589 12278 4292 12280
rect 2589 12275 2655 12278
rect 4286 12276 4292 12278
rect 4356 12338 4362 12340
rect 4981 12338 5047 12341
rect 4356 12336 5047 12338
rect 4356 12280 4986 12336
rect 5042 12280 5047 12336
rect 4356 12278 5047 12280
rect 4356 12276 4362 12278
rect 4981 12275 5047 12278
rect 6177 12336 6243 12341
rect 6177 12280 6182 12336
rect 6238 12280 6243 12336
rect 6177 12275 6243 12280
rect 6453 12338 6519 12341
rect 7557 12338 7623 12341
rect 6453 12336 7623 12338
rect 6453 12280 6458 12336
rect 6514 12280 7562 12336
rect 7618 12280 7623 12336
rect 6453 12278 7623 12280
rect 6453 12275 6519 12278
rect 7557 12275 7623 12278
rect 1710 12140 1716 12204
rect 1780 12202 1786 12204
rect 2405 12202 2471 12205
rect 1780 12200 2471 12202
rect 1780 12144 2410 12200
rect 2466 12144 2471 12200
rect 1780 12142 2471 12144
rect 1780 12140 1786 12142
rect 2405 12139 2471 12142
rect 3417 12202 3483 12205
rect 3734 12202 3740 12204
rect 3417 12200 3740 12202
rect 3417 12144 3422 12200
rect 3478 12144 3740 12200
rect 3417 12142 3740 12144
rect 3417 12139 3483 12142
rect 3734 12140 3740 12142
rect 3804 12140 3810 12204
rect 3877 12202 3943 12205
rect 4245 12202 4311 12205
rect 3877 12200 4311 12202
rect 3877 12144 3882 12200
rect 3938 12144 4250 12200
rect 4306 12144 4311 12200
rect 3877 12142 4311 12144
rect 3877 12139 3943 12142
rect 4245 12139 4311 12142
rect 4429 12202 4495 12205
rect 5073 12202 5139 12205
rect 4429 12200 5139 12202
rect 4429 12144 4434 12200
rect 4490 12144 5078 12200
rect 5134 12144 5139 12200
rect 4429 12142 5139 12144
rect 4429 12139 4495 12142
rect 5073 12139 5139 12142
rect 2313 12066 2379 12069
rect 3417 12066 3483 12069
rect 2313 12064 3483 12066
rect 2313 12008 2318 12064
rect 2374 12008 3422 12064
rect 3478 12008 3483 12064
rect 2313 12006 3483 12008
rect 2313 12003 2379 12006
rect 3417 12003 3483 12006
rect 3734 12004 3740 12068
rect 3804 12066 3810 12068
rect 4061 12066 4127 12069
rect 3804 12064 4127 12066
rect 3804 12008 4066 12064
rect 4122 12008 4127 12064
rect 3804 12006 4127 12008
rect 3804 12004 3810 12006
rect 4061 12003 4127 12006
rect 4286 12004 4292 12068
rect 4356 12066 4362 12068
rect 6180 12066 6240 12275
rect 6729 12204 6795 12205
rect 6678 12202 6684 12204
rect 6638 12142 6684 12202
rect 6748 12200 6795 12204
rect 6790 12144 6795 12200
rect 6678 12140 6684 12142
rect 6748 12140 6795 12144
rect 6729 12139 6795 12140
rect 6913 12202 6979 12205
rect 7744 12202 7804 12414
rect 8702 12412 8708 12414
rect 8772 12412 8778 12476
rect 9213 12474 9279 12477
rect 10688 12474 10748 12686
rect 12433 12683 12499 12686
rect 12893 12746 12959 12749
rect 13310 12746 13370 12822
rect 13813 12819 13879 12822
rect 14038 12820 14044 12884
rect 14108 12882 14114 12884
rect 14365 12882 14431 12885
rect 14108 12880 14431 12882
rect 14108 12824 14370 12880
rect 14426 12824 14431 12880
rect 14108 12822 14431 12824
rect 14108 12820 14114 12822
rect 14365 12819 14431 12822
rect 15469 12884 15535 12885
rect 15469 12880 15516 12884
rect 15580 12882 15586 12884
rect 15469 12824 15474 12880
rect 15469 12820 15516 12824
rect 15580 12822 15626 12882
rect 15580 12820 15586 12822
rect 15469 12819 15535 12820
rect 12893 12744 13370 12746
rect 12893 12688 12898 12744
rect 12954 12688 13370 12744
rect 12893 12686 13370 12688
rect 14181 12746 14247 12749
rect 14825 12746 14891 12749
rect 14181 12744 14891 12746
rect 14181 12688 14186 12744
rect 14242 12688 14830 12744
rect 14886 12688 14891 12744
rect 14181 12686 14891 12688
rect 12893 12683 12959 12686
rect 14181 12683 14247 12686
rect 14825 12683 14891 12686
rect 11513 12610 11579 12613
rect 13997 12610 14063 12613
rect 11513 12608 13738 12610
rect 11513 12552 11518 12608
rect 11574 12552 13738 12608
rect 11513 12550 13738 12552
rect 11513 12547 11579 12550
rect 10816 12544 11132 12545
rect 10816 12480 10822 12544
rect 10886 12480 10902 12544
rect 10966 12480 10982 12544
rect 11046 12480 11062 12544
rect 11126 12480 11132 12544
rect 10816 12479 11132 12480
rect 9213 12472 10748 12474
rect 9213 12416 9218 12472
rect 9274 12416 10748 12472
rect 9213 12414 10748 12416
rect 9213 12411 9279 12414
rect 11462 12412 11468 12476
rect 11532 12474 11538 12476
rect 11789 12474 11855 12477
rect 11532 12472 11855 12474
rect 11532 12416 11794 12472
rect 11850 12416 11855 12472
rect 11532 12414 11855 12416
rect 11532 12412 11538 12414
rect 11789 12411 11855 12414
rect 12249 12474 12315 12477
rect 13169 12474 13235 12477
rect 12249 12472 13235 12474
rect 12249 12416 12254 12472
rect 12310 12416 13174 12472
rect 13230 12416 13235 12472
rect 12249 12414 13235 12416
rect 12249 12411 12315 12414
rect 13169 12411 13235 12414
rect 13678 12440 13738 12550
rect 13862 12608 14063 12610
rect 13862 12552 14002 12608
rect 14058 12552 14063 12608
rect 13862 12550 14063 12552
rect 13862 12440 13922 12550
rect 13997 12547 14063 12550
rect 15377 12610 15443 12613
rect 15510 12610 15516 12612
rect 15377 12608 15516 12610
rect 15377 12552 15382 12608
rect 15438 12552 15516 12608
rect 15377 12550 15516 12552
rect 15377 12547 15443 12550
rect 15510 12548 15516 12550
rect 15580 12548 15586 12612
rect 14764 12544 15080 12545
rect 14764 12480 14770 12544
rect 14834 12480 14850 12544
rect 14914 12480 14930 12544
rect 14994 12480 15010 12544
rect 15074 12480 15080 12544
rect 14764 12479 15080 12480
rect 13678 12380 13922 12440
rect 9581 12336 9647 12341
rect 9581 12280 9586 12336
rect 9642 12280 9647 12336
rect 9581 12275 9647 12280
rect 9765 12338 9831 12341
rect 10133 12338 10199 12341
rect 9765 12336 10199 12338
rect 9765 12280 9770 12336
rect 9826 12280 10138 12336
rect 10194 12280 10199 12336
rect 9765 12278 10199 12280
rect 9765 12275 9831 12278
rect 10133 12275 10199 12278
rect 10358 12276 10364 12340
rect 10428 12338 10434 12340
rect 11053 12338 11119 12341
rect 11462 12338 11468 12340
rect 10428 12278 10978 12338
rect 10428 12276 10434 12278
rect 9584 12205 9644 12275
rect 6913 12200 7804 12202
rect 6913 12144 6918 12200
rect 6974 12144 7804 12200
rect 6913 12142 7804 12144
rect 6913 12139 6979 12142
rect 7966 12140 7972 12204
rect 8036 12202 8042 12204
rect 8201 12202 8267 12205
rect 8036 12200 8267 12202
rect 8036 12144 8206 12200
rect 8262 12144 8267 12200
rect 8036 12142 8267 12144
rect 8036 12140 8042 12142
rect 8201 12139 8267 12142
rect 8569 12202 8635 12205
rect 9029 12202 9095 12205
rect 8569 12200 9095 12202
rect 8569 12144 8574 12200
rect 8630 12144 9034 12200
rect 9090 12144 9095 12200
rect 8569 12142 9095 12144
rect 8569 12139 8635 12142
rect 9029 12139 9095 12142
rect 9581 12200 9647 12205
rect 9581 12144 9586 12200
rect 9642 12144 9647 12200
rect 9581 12139 9647 12144
rect 9765 12204 9831 12205
rect 9765 12200 9812 12204
rect 9876 12202 9882 12204
rect 10918 12202 10978 12278
rect 11053 12336 11468 12338
rect 11053 12280 11058 12336
rect 11114 12280 11468 12336
rect 11053 12278 11468 12280
rect 11053 12275 11119 12278
rect 11462 12276 11468 12278
rect 11532 12276 11538 12340
rect 13445 12338 13511 12341
rect 11654 12336 13511 12338
rect 11654 12280 13450 12336
rect 13506 12280 13511 12336
rect 11654 12278 13511 12280
rect 11654 12202 11714 12278
rect 13445 12275 13511 12278
rect 14089 12338 14155 12341
rect 14089 12336 14428 12338
rect 14089 12280 14094 12336
rect 14150 12280 14428 12336
rect 14089 12278 14428 12280
rect 14089 12275 14155 12278
rect 14368 12205 14428 12278
rect 14038 12202 14044 12204
rect 9765 12144 9770 12200
rect 9765 12140 9812 12144
rect 9876 12142 10794 12202
rect 10918 12142 11714 12202
rect 11792 12142 14044 12202
rect 9876 12140 9882 12142
rect 9765 12139 9831 12140
rect 8702 12066 8708 12068
rect 4356 12006 4492 12066
rect 6180 12006 8708 12066
rect 4356 12004 4362 12006
rect 2589 11932 2655 11933
rect 2589 11928 2636 11932
rect 2700 11930 2706 11932
rect 3141 11930 3207 11933
rect 4286 11930 4292 11932
rect 2589 11872 2594 11928
rect 2589 11868 2636 11872
rect 2700 11870 2746 11930
rect 3141 11928 4292 11930
rect 3141 11872 3146 11928
rect 3202 11872 4292 11928
rect 3141 11870 4292 11872
rect 2700 11868 2706 11870
rect 2589 11867 2655 11868
rect 3141 11867 3207 11870
rect 4286 11868 4292 11870
rect 4356 11868 4362 11932
rect 2221 11796 2287 11797
rect 2221 11792 2268 11796
rect 2332 11794 2338 11796
rect 4061 11794 4127 11797
rect 4432 11794 4492 12006
rect 8702 12004 8708 12006
rect 8772 12004 8778 12068
rect 9397 12066 9463 12069
rect 9581 12066 9647 12069
rect 9397 12064 9647 12066
rect 9397 12008 9402 12064
rect 9458 12008 9586 12064
rect 9642 12008 9647 12064
rect 9397 12006 9647 12008
rect 9397 12003 9463 12006
rect 9581 12003 9647 12006
rect 9806 12004 9812 12068
rect 9876 12066 9882 12068
rect 10225 12066 10291 12069
rect 9876 12064 10291 12066
rect 9876 12008 10230 12064
rect 10286 12008 10291 12064
rect 9876 12006 10291 12008
rect 9876 12004 9882 12006
rect 10225 12003 10291 12006
rect 10358 12004 10364 12068
rect 10428 12066 10434 12068
rect 10593 12066 10659 12069
rect 10428 12064 10659 12066
rect 10428 12008 10598 12064
rect 10654 12008 10659 12064
rect 10428 12006 10659 12008
rect 10734 12066 10794 12142
rect 11792 12066 11852 12142
rect 14038 12140 14044 12142
rect 14108 12140 14114 12204
rect 14365 12200 14431 12205
rect 14365 12144 14370 12200
rect 14426 12144 14431 12200
rect 14365 12139 14431 12144
rect 14733 12202 14799 12205
rect 15142 12202 15148 12204
rect 14733 12200 15148 12202
rect 14733 12144 14738 12200
rect 14794 12144 15148 12200
rect 14733 12142 15148 12144
rect 14733 12139 14799 12142
rect 15142 12140 15148 12142
rect 15212 12140 15218 12204
rect 15653 12202 15719 12205
rect 16246 12202 16252 12204
rect 15653 12200 16252 12202
rect 15653 12144 15658 12200
rect 15714 12144 16252 12200
rect 15653 12142 16252 12144
rect 15653 12139 15719 12142
rect 16246 12140 16252 12142
rect 16316 12140 16322 12204
rect 10734 12006 11852 12066
rect 12249 12066 12315 12069
rect 12382 12066 12388 12068
rect 12249 12064 12388 12066
rect 12249 12008 12254 12064
rect 12310 12008 12388 12064
rect 12249 12006 12388 12008
rect 10428 12004 10434 12006
rect 10593 12003 10659 12006
rect 12249 12003 12315 12006
rect 12382 12004 12388 12006
rect 12452 12004 12458 12068
rect 13721 12066 13787 12069
rect 13310 12064 13787 12066
rect 13310 12008 13726 12064
rect 13782 12008 13787 12064
rect 13310 12006 13787 12008
rect 4894 12000 5210 12001
rect 4894 11936 4900 12000
rect 4964 11936 4980 12000
rect 5044 11936 5060 12000
rect 5124 11936 5140 12000
rect 5204 11936 5210 12000
rect 4894 11935 5210 11936
rect 8842 12000 9158 12001
rect 8842 11936 8848 12000
rect 8912 11936 8928 12000
rect 8992 11936 9008 12000
rect 9072 11936 9088 12000
rect 9152 11936 9158 12000
rect 8842 11935 9158 11936
rect 12790 12000 13106 12001
rect 12790 11936 12796 12000
rect 12860 11936 12876 12000
rect 12940 11936 12956 12000
rect 13020 11936 13036 12000
rect 13100 11936 13106 12000
rect 12790 11935 13106 11936
rect 5993 11930 6059 11933
rect 7276 11930 7282 11932
rect 5993 11928 7282 11930
rect 5993 11872 5998 11928
rect 6054 11872 7282 11928
rect 5993 11870 7282 11872
rect 5993 11867 6059 11870
rect 7276 11868 7282 11870
rect 7346 11868 7352 11932
rect 10225 11930 10291 11933
rect 10961 11930 11027 11933
rect 10225 11928 11027 11930
rect 10225 11872 10230 11928
rect 10286 11872 10966 11928
rect 11022 11872 11027 11928
rect 10225 11870 11027 11872
rect 10225 11867 10291 11870
rect 10961 11867 11027 11870
rect 11697 11930 11763 11933
rect 12341 11932 12407 11933
rect 11697 11928 12266 11930
rect 11697 11872 11702 11928
rect 11758 11872 12266 11928
rect 11697 11870 12266 11872
rect 11697 11867 11763 11870
rect 2221 11736 2226 11792
rect 2221 11732 2268 11736
rect 2332 11734 2378 11794
rect 4061 11792 4492 11794
rect 4061 11736 4066 11792
rect 4122 11736 4492 11792
rect 4061 11734 4492 11736
rect 5165 11794 5231 11797
rect 5390 11794 5396 11796
rect 5165 11792 5396 11794
rect 5165 11736 5170 11792
rect 5226 11736 5396 11792
rect 5165 11734 5396 11736
rect 2332 11732 2338 11734
rect 2221 11731 2287 11732
rect 4061 11731 4127 11734
rect 5165 11731 5231 11734
rect 5390 11732 5396 11734
rect 5460 11732 5466 11796
rect 6637 11794 6703 11797
rect 12065 11794 12131 11797
rect 6637 11792 12131 11794
rect 6637 11736 6642 11792
rect 6698 11736 12070 11792
rect 12126 11736 12131 11792
rect 6637 11734 12131 11736
rect 12206 11794 12266 11870
rect 12341 11928 12388 11932
rect 12452 11930 12458 11932
rect 12341 11872 12346 11928
rect 12341 11868 12388 11872
rect 12452 11870 12498 11930
rect 12452 11868 12458 11870
rect 12341 11867 12407 11868
rect 13310 11794 13370 12006
rect 13721 12003 13787 12006
rect 14038 12004 14044 12068
rect 14108 12066 14114 12068
rect 14917 12066 14983 12069
rect 14108 12064 14983 12066
rect 14108 12008 14922 12064
rect 14978 12008 14983 12064
rect 14108 12006 14983 12008
rect 14108 12004 14114 12006
rect 14917 12003 14983 12006
rect 13445 11930 13511 11933
rect 14825 11930 14891 11933
rect 13445 11928 14891 11930
rect 13445 11872 13450 11928
rect 13506 11872 14830 11928
rect 14886 11872 14891 11928
rect 13445 11870 14891 11872
rect 13445 11867 13511 11870
rect 14825 11867 14891 11870
rect 12206 11734 13370 11794
rect 6637 11731 6703 11734
rect 12065 11731 12131 11734
rect 13854 11732 13860 11796
rect 13924 11794 13930 11796
rect 15142 11794 15148 11796
rect 13924 11734 15148 11794
rect 13924 11732 13930 11734
rect 15142 11732 15148 11734
rect 15212 11732 15218 11796
rect 8518 11658 8524 11660
rect 2730 11598 8524 11658
rect 0 11250 400 11280
rect 2730 11250 2790 11598
rect 8518 11596 8524 11598
rect 8588 11596 8594 11660
rect 8702 11596 8708 11660
rect 8772 11658 8778 11660
rect 10869 11658 10935 11661
rect 8772 11656 10935 11658
rect 8772 11600 10874 11656
rect 10930 11600 10935 11656
rect 8772 11598 10935 11600
rect 8772 11596 8778 11598
rect 10869 11595 10935 11598
rect 11053 11658 11119 11661
rect 13854 11658 13860 11660
rect 11053 11656 13860 11658
rect 11053 11600 11058 11656
rect 11114 11600 13860 11656
rect 11053 11598 13860 11600
rect 11053 11595 11119 11598
rect 13854 11596 13860 11598
rect 13924 11596 13930 11660
rect 15694 11658 15700 11660
rect 14230 11598 15700 11658
rect 4153 11522 4219 11525
rect 5073 11522 5139 11525
rect 6310 11522 6316 11524
rect 4153 11520 6316 11522
rect 4153 11464 4158 11520
rect 4214 11464 5078 11520
rect 5134 11464 6316 11520
rect 4153 11462 6316 11464
rect 4153 11459 4219 11462
rect 5073 11459 5139 11462
rect 6310 11460 6316 11462
rect 6380 11460 6386 11524
rect 8150 11460 8156 11524
rect 8220 11522 8226 11524
rect 8518 11522 8524 11524
rect 8220 11462 8524 11522
rect 8220 11460 8226 11462
rect 8518 11460 8524 11462
rect 8588 11460 8594 11524
rect 11697 11522 11763 11525
rect 11830 11522 11836 11524
rect 11697 11520 11836 11522
rect 11697 11464 11702 11520
rect 11758 11464 11836 11520
rect 11697 11462 11836 11464
rect 11697 11459 11763 11462
rect 11830 11460 11836 11462
rect 11900 11460 11906 11524
rect 13164 11522 13170 11524
rect 12252 11462 13170 11522
rect 2920 11456 3236 11457
rect 2920 11392 2926 11456
rect 2990 11392 3006 11456
rect 3070 11392 3086 11456
rect 3150 11392 3166 11456
rect 3230 11392 3236 11456
rect 2920 11391 3236 11392
rect 6868 11456 7184 11457
rect 6868 11392 6874 11456
rect 6938 11392 6954 11456
rect 7018 11392 7034 11456
rect 7098 11392 7114 11456
rect 7178 11392 7184 11456
rect 6868 11391 7184 11392
rect 10816 11456 11132 11457
rect 10816 11392 10822 11456
rect 10886 11392 10902 11456
rect 10966 11392 10982 11456
rect 11046 11392 11062 11456
rect 11126 11392 11132 11456
rect 10816 11391 11132 11392
rect 12252 11389 12312 11462
rect 13164 11460 13170 11462
rect 13234 11460 13240 11524
rect 13721 11522 13787 11525
rect 14038 11522 14044 11524
rect 13721 11520 14044 11522
rect 13721 11464 13726 11520
rect 13782 11464 14044 11520
rect 13721 11462 14044 11464
rect 13721 11459 13787 11462
rect 14038 11460 14044 11462
rect 14108 11460 14114 11524
rect 3366 11324 3372 11388
rect 3436 11386 3442 11388
rect 3601 11386 3667 11389
rect 3436 11384 3667 11386
rect 3436 11328 3606 11384
rect 3662 11328 3667 11384
rect 3436 11326 3667 11328
rect 3436 11324 3442 11326
rect 3601 11323 3667 11326
rect 4061 11386 4127 11389
rect 4061 11384 4584 11386
rect 4061 11328 4066 11384
rect 4122 11328 4584 11384
rect 4061 11326 4584 11328
rect 4061 11323 4127 11326
rect 0 11190 2790 11250
rect 2957 11250 3023 11253
rect 3550 11250 3556 11252
rect 2957 11248 3556 11250
rect 2957 11192 2962 11248
rect 3018 11192 3556 11248
rect 2957 11190 3556 11192
rect 0 11160 400 11190
rect 2957 11187 3023 11190
rect 3550 11188 3556 11190
rect 3620 11250 3626 11252
rect 4245 11250 4311 11253
rect 3620 11248 4311 11250
rect 3620 11192 4250 11248
rect 4306 11192 4311 11248
rect 3620 11190 4311 11192
rect 4524 11250 4584 11326
rect 4654 11324 4660 11388
rect 4724 11386 4730 11388
rect 4797 11386 4863 11389
rect 4724 11384 4863 11386
rect 4724 11328 4802 11384
rect 4858 11328 4863 11384
rect 4724 11326 4863 11328
rect 4724 11324 4730 11326
rect 4797 11323 4863 11326
rect 7373 11384 7439 11389
rect 7373 11328 7378 11384
rect 7434 11328 7439 11384
rect 7373 11323 7439 11328
rect 8201 11386 8267 11389
rect 9254 11386 9260 11388
rect 8201 11384 9260 11386
rect 8201 11328 8206 11384
rect 8262 11328 9260 11384
rect 8201 11326 9260 11328
rect 8201 11323 8267 11326
rect 9254 11324 9260 11326
rect 9324 11324 9330 11388
rect 12249 11384 12315 11389
rect 12249 11328 12254 11384
rect 12310 11328 12315 11384
rect 12249 11323 12315 11328
rect 12525 11386 12591 11389
rect 14230 11386 14290 11598
rect 15694 11596 15700 11598
rect 15764 11596 15770 11660
rect 14764 11456 15080 11457
rect 14764 11392 14770 11456
rect 14834 11392 14850 11456
rect 14914 11392 14930 11456
rect 14994 11392 15010 11456
rect 15074 11392 15080 11456
rect 14764 11391 15080 11392
rect 12525 11384 14290 11386
rect 12525 11328 12530 11384
rect 12586 11328 14290 11384
rect 12525 11326 14290 11328
rect 12525 11323 12591 11326
rect 5942 11250 5948 11252
rect 4524 11190 5948 11250
rect 3620 11188 3626 11190
rect 4245 11187 4311 11190
rect 5942 11188 5948 11190
rect 6012 11250 6018 11252
rect 7097 11250 7163 11253
rect 6012 11248 7163 11250
rect 6012 11192 7102 11248
rect 7158 11192 7163 11248
rect 6012 11190 7163 11192
rect 7376 11250 7436 11323
rect 8150 11250 8156 11252
rect 7376 11190 8156 11250
rect 6012 11188 6018 11190
rect 7097 11187 7163 11190
rect 8150 11188 8156 11190
rect 8220 11188 8226 11252
rect 9305 11250 9371 11253
rect 8296 11248 9371 11250
rect 8296 11192 9310 11248
rect 9366 11192 9371 11248
rect 8296 11190 9371 11192
rect 2446 11052 2452 11116
rect 2516 11114 2522 11116
rect 2865 11114 2931 11117
rect 8296 11114 8356 11190
rect 9305 11187 9371 11190
rect 9581 11250 9647 11253
rect 11421 11250 11487 11253
rect 15285 11250 15351 11253
rect 9581 11248 11487 11250
rect 9581 11192 9586 11248
rect 9642 11192 11426 11248
rect 11482 11192 11487 11248
rect 12436 11248 15351 11250
rect 12436 11216 15290 11248
rect 9581 11190 11487 11192
rect 9581 11187 9647 11190
rect 11421 11187 11487 11190
rect 12344 11192 15290 11216
rect 15346 11192 15351 11248
rect 12344 11190 15351 11192
rect 12344 11156 12496 11190
rect 15285 11187 15351 11190
rect 2516 11112 2931 11114
rect 2516 11056 2870 11112
rect 2926 11056 2931 11112
rect 2516 11054 2931 11056
rect 2516 11052 2522 11054
rect 2865 11051 2931 11054
rect 3006 11054 8356 11114
rect 9029 11114 9095 11117
rect 10593 11114 10659 11117
rect 9029 11112 10659 11114
rect 9029 11056 9034 11112
rect 9090 11056 10598 11112
rect 10654 11056 10659 11112
rect 9029 11054 10659 11056
rect 2589 10842 2655 10845
rect 3006 10842 3066 11054
rect 9029 11051 9095 11054
rect 10593 11051 10659 11054
rect 11462 11052 11468 11116
rect 11532 11114 11538 11116
rect 12157 11114 12223 11117
rect 11532 11112 12223 11114
rect 11532 11056 12162 11112
rect 12218 11056 12223 11112
rect 11532 11054 12223 11056
rect 11532 11052 11538 11054
rect 12157 11051 12223 11054
rect 3877 10980 3943 10981
rect 4705 10980 4771 10981
rect 3877 10976 3924 10980
rect 3988 10978 3994 10980
rect 3877 10920 3882 10976
rect 3877 10916 3924 10920
rect 3988 10918 4034 10978
rect 3988 10916 3994 10918
rect 4654 10916 4660 10980
rect 4724 10978 4771 10980
rect 8477 10978 8543 10981
rect 8702 10978 8708 10980
rect 4724 10976 4816 10978
rect 4766 10920 4816 10976
rect 4724 10918 4816 10920
rect 8477 10976 8708 10978
rect 8477 10920 8482 10976
rect 8538 10920 8708 10976
rect 8477 10918 8708 10920
rect 4724 10916 4771 10918
rect 3877 10915 3943 10916
rect 4705 10915 4771 10916
rect 8477 10915 8543 10918
rect 8702 10916 8708 10918
rect 8772 10916 8778 10980
rect 9673 10978 9739 10981
rect 10174 10978 10180 10980
rect 9673 10976 10180 10978
rect 9673 10920 9678 10976
rect 9734 10920 10180 10976
rect 9673 10918 10180 10920
rect 9673 10915 9739 10918
rect 10174 10916 10180 10918
rect 10244 10916 10250 10980
rect 10961 10978 11027 10981
rect 11462 10978 11468 10980
rect 10961 10976 11468 10978
rect 10961 10920 10966 10976
rect 11022 10920 11468 10976
rect 10961 10918 11468 10920
rect 10961 10915 11027 10918
rect 11462 10916 11468 10918
rect 11532 10916 11538 10980
rect 12344 10978 12404 11156
rect 14406 11114 14412 11116
rect 11838 10918 12404 10978
rect 12574 11054 14412 11114
rect 4894 10912 5210 10913
rect 4894 10848 4900 10912
rect 4964 10848 4980 10912
rect 5044 10848 5060 10912
rect 5124 10848 5140 10912
rect 5204 10848 5210 10912
rect 4894 10847 5210 10848
rect 8842 10912 9158 10913
rect 8842 10848 8848 10912
rect 8912 10848 8928 10912
rect 8992 10848 9008 10912
rect 9072 10848 9088 10912
rect 9152 10848 9158 10912
rect 8842 10847 9158 10848
rect 2589 10840 3066 10842
rect 2589 10784 2594 10840
rect 2650 10784 3066 10840
rect 2589 10782 3066 10784
rect 10593 10842 10659 10845
rect 11838 10844 11898 10918
rect 11830 10842 11836 10844
rect 10593 10840 11836 10842
rect 10593 10784 10598 10840
rect 10654 10784 11836 10840
rect 10593 10782 11836 10784
rect 2589 10779 2655 10782
rect 10593 10779 10659 10782
rect 11830 10780 11836 10782
rect 11900 10780 11906 10844
rect 12249 10842 12315 10845
rect 12574 10842 12634 11054
rect 14406 11052 14412 11054
rect 14476 11052 14482 11116
rect 14917 11114 14983 11117
rect 15878 11114 15884 11116
rect 14917 11112 15884 11114
rect 14917 11056 14922 11112
rect 14978 11056 15884 11112
rect 14917 11054 15884 11056
rect 14917 11051 14983 11054
rect 15878 11052 15884 11054
rect 15948 11052 15954 11116
rect 13261 10978 13327 10981
rect 13997 10978 14063 10981
rect 13261 10976 14063 10978
rect 13261 10920 13266 10976
rect 13322 10920 14002 10976
rect 14058 10920 14063 10976
rect 13261 10918 14063 10920
rect 13261 10915 13327 10918
rect 13997 10915 14063 10918
rect 14641 10978 14707 10981
rect 15193 10978 15259 10981
rect 14641 10976 15259 10978
rect 14641 10920 14646 10976
rect 14702 10920 15198 10976
rect 15254 10920 15259 10976
rect 14641 10918 15259 10920
rect 14641 10915 14707 10918
rect 15193 10915 15259 10918
rect 12790 10912 13106 10913
rect 12790 10848 12796 10912
rect 12860 10848 12876 10912
rect 12940 10848 12956 10912
rect 13020 10848 13036 10912
rect 13100 10848 13106 10912
rect 12790 10847 13106 10848
rect 12249 10840 12634 10842
rect 12249 10784 12254 10840
rect 12310 10784 12634 10840
rect 12249 10782 12634 10784
rect 12249 10779 12315 10782
rect 14038 10780 14044 10844
rect 14108 10842 14114 10844
rect 14825 10842 14891 10845
rect 14108 10840 14891 10842
rect 14108 10784 14830 10840
rect 14886 10784 14891 10840
rect 14108 10782 14891 10784
rect 14108 10780 14114 10782
rect 14825 10779 14891 10782
rect 15285 10842 15351 10845
rect 15694 10842 15700 10844
rect 15285 10840 15700 10842
rect 15285 10784 15290 10840
rect 15346 10784 15700 10840
rect 15285 10782 15700 10784
rect 15285 10779 15351 10782
rect 15694 10780 15700 10782
rect 15764 10780 15770 10844
rect 1761 10706 1827 10709
rect 1894 10706 1900 10708
rect 1761 10704 1900 10706
rect 1761 10648 1766 10704
rect 1822 10648 1900 10704
rect 1761 10646 1900 10648
rect 1761 10643 1827 10646
rect 1894 10644 1900 10646
rect 1964 10644 1970 10708
rect 4429 10706 4495 10709
rect 8385 10706 8451 10709
rect 4429 10704 8451 10706
rect 4429 10648 4434 10704
rect 4490 10648 8390 10704
rect 8446 10648 8451 10704
rect 4429 10646 8451 10648
rect 4429 10643 4495 10646
rect 8385 10643 8451 10646
rect 9029 10706 9095 10709
rect 9438 10706 9444 10708
rect 9029 10704 9444 10706
rect 9029 10648 9034 10704
rect 9090 10648 9444 10704
rect 9029 10646 9444 10648
rect 9029 10643 9095 10646
rect 9438 10644 9444 10646
rect 9508 10644 9514 10708
rect 9990 10644 9996 10708
rect 10060 10706 10066 10708
rect 10133 10706 10199 10709
rect 10060 10704 10199 10706
rect 10060 10648 10138 10704
rect 10194 10648 10199 10704
rect 10060 10646 10199 10648
rect 10060 10644 10066 10646
rect 10133 10643 10199 10646
rect 10358 10644 10364 10708
rect 10428 10706 10434 10708
rect 15009 10706 15075 10709
rect 15469 10706 15535 10709
rect 10428 10704 15535 10706
rect 10428 10648 15014 10704
rect 15070 10648 15474 10704
rect 15530 10648 15535 10704
rect 10428 10646 15535 10648
rect 10428 10644 10434 10646
rect 15009 10643 15075 10646
rect 15469 10643 15535 10646
rect 2221 10570 2287 10573
rect 4705 10570 4771 10573
rect 2221 10568 4771 10570
rect 2221 10512 2226 10568
rect 2282 10512 4710 10568
rect 4766 10512 4771 10568
rect 2221 10510 4771 10512
rect 2221 10507 2287 10510
rect 4705 10507 4771 10510
rect 4889 10570 4955 10573
rect 5574 10570 5580 10572
rect 4889 10568 5580 10570
rect 4889 10512 4894 10568
rect 4950 10512 5580 10568
rect 4889 10510 5580 10512
rect 4889 10507 4955 10510
rect 5574 10508 5580 10510
rect 5644 10508 5650 10572
rect 6126 10508 6132 10572
rect 6196 10570 6202 10572
rect 6196 10510 7712 10570
rect 6196 10508 6202 10510
rect 3509 10434 3575 10437
rect 3374 10432 3575 10434
rect 3374 10376 3514 10432
rect 3570 10376 3575 10432
rect 3374 10374 3575 10376
rect 2920 10368 3236 10369
rect 2920 10304 2926 10368
rect 2990 10304 3006 10368
rect 3070 10304 3086 10368
rect 3150 10304 3166 10368
rect 3230 10304 3236 10368
rect 2920 10303 3236 10304
rect 3141 10162 3207 10165
rect 3374 10162 3434 10374
rect 3509 10371 3575 10374
rect 4102 10372 4108 10436
rect 4172 10434 4178 10436
rect 6177 10434 6243 10437
rect 4172 10432 6243 10434
rect 4172 10376 6182 10432
rect 6238 10376 6243 10432
rect 4172 10374 6243 10376
rect 7652 10434 7712 10510
rect 7782 10508 7788 10572
rect 7852 10570 7858 10572
rect 7852 10510 11944 10570
rect 7852 10508 7858 10510
rect 9438 10434 9444 10436
rect 7652 10374 9444 10434
rect 4172 10372 4178 10374
rect 6177 10371 6243 10374
rect 9438 10372 9444 10374
rect 9508 10372 9514 10436
rect 9765 10434 9831 10437
rect 10174 10434 10180 10436
rect 9765 10432 10180 10434
rect 9765 10376 9770 10432
rect 9826 10376 10180 10432
rect 9765 10374 10180 10376
rect 9765 10371 9831 10374
rect 10174 10372 10180 10374
rect 10244 10372 10250 10436
rect 11329 10434 11395 10437
rect 11462 10434 11468 10436
rect 11329 10432 11468 10434
rect 11329 10376 11334 10432
rect 11390 10376 11468 10432
rect 11329 10374 11468 10376
rect 11329 10371 11395 10374
rect 11462 10372 11468 10374
rect 11532 10372 11538 10436
rect 11884 10434 11944 10510
rect 12014 10508 12020 10572
rect 12084 10570 12090 10572
rect 12801 10570 12867 10573
rect 12084 10568 12867 10570
rect 12084 10512 12806 10568
rect 12862 10512 12867 10568
rect 12084 10510 12867 10512
rect 12084 10508 12090 10510
rect 12801 10507 12867 10510
rect 13169 10570 13235 10573
rect 14733 10570 14799 10573
rect 13169 10568 14799 10570
rect 13169 10512 13174 10568
rect 13230 10512 14738 10568
rect 14794 10512 14799 10568
rect 13169 10510 14799 10512
rect 13169 10507 13235 10510
rect 14733 10507 14799 10510
rect 13353 10434 13419 10437
rect 11884 10432 13419 10434
rect 11884 10376 13358 10432
rect 13414 10376 13419 10432
rect 11884 10374 13419 10376
rect 13353 10371 13419 10374
rect 13905 10432 13971 10437
rect 13905 10376 13910 10432
rect 13966 10376 13971 10432
rect 13905 10371 13971 10376
rect 14273 10434 14339 10437
rect 14590 10434 14596 10436
rect 14273 10432 14596 10434
rect 14273 10376 14278 10432
rect 14334 10376 14596 10432
rect 14273 10374 14596 10376
rect 14273 10371 14339 10374
rect 14590 10372 14596 10374
rect 14660 10372 14666 10436
rect 15653 10434 15719 10437
rect 15288 10432 15719 10434
rect 15288 10376 15658 10432
rect 15714 10376 15719 10432
rect 15288 10374 15719 10376
rect 6868 10368 7184 10369
rect 6868 10304 6874 10368
rect 6938 10304 6954 10368
rect 7018 10304 7034 10368
rect 7098 10304 7114 10368
rect 7178 10304 7184 10368
rect 6868 10303 7184 10304
rect 10816 10368 11132 10369
rect 10816 10304 10822 10368
rect 10886 10304 10902 10368
rect 10966 10304 10982 10368
rect 11046 10304 11062 10368
rect 11126 10304 11132 10368
rect 10816 10303 11132 10304
rect 4613 10298 4679 10301
rect 5993 10298 6059 10301
rect 4613 10296 6059 10298
rect 4613 10240 4618 10296
rect 4674 10240 5998 10296
rect 6054 10240 6059 10296
rect 4613 10238 6059 10240
rect 4613 10235 4679 10238
rect 5993 10235 6059 10238
rect 8293 10296 8359 10301
rect 8293 10240 8298 10296
rect 8354 10240 8359 10296
rect 8293 10235 8359 10240
rect 11237 10298 11303 10301
rect 13445 10298 13511 10301
rect 11237 10296 13511 10298
rect 11237 10240 11242 10296
rect 11298 10240 13450 10296
rect 13506 10240 13511 10296
rect 11237 10238 13511 10240
rect 13908 10298 13968 10371
rect 14764 10368 15080 10369
rect 14764 10304 14770 10368
rect 14834 10304 14850 10368
rect 14914 10304 14930 10368
rect 14994 10304 15010 10368
rect 15074 10304 15080 10368
rect 14764 10303 15080 10304
rect 15288 10301 15348 10374
rect 15653 10371 15719 10374
rect 13908 10238 14704 10298
rect 11237 10235 11303 10238
rect 13445 10235 13511 10238
rect 3141 10160 3434 10162
rect 3141 10104 3146 10160
rect 3202 10104 3434 10160
rect 3141 10102 3434 10104
rect 3141 10099 3207 10102
rect 4286 10100 4292 10164
rect 4356 10162 4362 10164
rect 5993 10162 6059 10165
rect 4356 10160 6059 10162
rect 4356 10104 5998 10160
rect 6054 10104 6059 10160
rect 4356 10102 6059 10104
rect 4356 10100 4362 10102
rect 5993 10099 6059 10102
rect 3141 10026 3207 10029
rect 5717 10026 5783 10029
rect 8109 10026 8175 10029
rect 3141 10024 8175 10026
rect 3141 9968 3146 10024
rect 3202 9968 5722 10024
rect 5778 9968 8114 10024
rect 8170 9968 8175 10024
rect 3141 9966 8175 9968
rect 3141 9963 3207 9966
rect 5717 9963 5783 9966
rect 8109 9963 8175 9966
rect 6126 9828 6132 9892
rect 6196 9890 6202 9892
rect 8296 9890 8356 10235
rect 8518 10100 8524 10164
rect 8588 10162 8594 10164
rect 14181 10162 14247 10165
rect 8588 10160 14247 10162
rect 8588 10104 14186 10160
rect 14242 10104 14247 10160
rect 8588 10102 14247 10104
rect 14644 10162 14704 10238
rect 15285 10296 15351 10301
rect 15285 10240 15290 10296
rect 15346 10240 15351 10296
rect 15285 10235 15351 10240
rect 15561 10162 15627 10165
rect 14644 10160 15627 10162
rect 14644 10104 15566 10160
rect 15622 10104 15627 10160
rect 14644 10102 15627 10104
rect 8588 10100 8594 10102
rect 14181 10099 14247 10102
rect 15561 10099 15627 10102
rect 9213 10026 9279 10029
rect 9213 10024 9920 10026
rect 9213 9968 9218 10024
rect 9274 9968 9920 10024
rect 9213 9966 9920 9968
rect 9213 9963 9279 9966
rect 8569 9890 8635 9893
rect 6196 9888 8635 9890
rect 6196 9832 8574 9888
rect 8630 9832 8635 9888
rect 6196 9830 8635 9832
rect 9860 9890 9920 9966
rect 9990 9964 9996 10028
rect 10060 10026 10066 10028
rect 12985 10026 13051 10029
rect 15101 10026 15167 10029
rect 10060 10024 15167 10026
rect 10060 9968 12990 10024
rect 13046 9968 15106 10024
rect 15162 9968 15167 10024
rect 10060 9966 15167 9968
rect 10060 9964 10066 9966
rect 12985 9963 13051 9966
rect 15101 9963 15167 9966
rect 12525 9890 12591 9893
rect 9860 9888 12591 9890
rect 9860 9832 12530 9888
rect 12586 9832 12591 9888
rect 9860 9830 12591 9832
rect 6196 9828 6202 9830
rect 8569 9827 8635 9830
rect 12525 9827 12591 9830
rect 13445 9890 13511 9893
rect 14089 9890 14155 9893
rect 13445 9888 14155 9890
rect 13445 9832 13450 9888
rect 13506 9832 14094 9888
rect 14150 9832 14155 9888
rect 13445 9830 14155 9832
rect 13445 9827 13511 9830
rect 14089 9827 14155 9830
rect 14273 9890 14339 9893
rect 14549 9890 14615 9893
rect 14273 9888 14615 9890
rect 14273 9832 14278 9888
rect 14334 9832 14554 9888
rect 14610 9832 14615 9888
rect 14273 9830 14615 9832
rect 14273 9827 14339 9830
rect 14549 9827 14615 9830
rect 14825 9890 14891 9893
rect 16430 9890 16436 9892
rect 14825 9888 16436 9890
rect 14825 9832 14830 9888
rect 14886 9832 16436 9888
rect 14825 9830 16436 9832
rect 14825 9827 14891 9830
rect 16430 9828 16436 9830
rect 16500 9828 16506 9892
rect 4894 9824 5210 9825
rect 0 9754 400 9784
rect 4894 9760 4900 9824
rect 4964 9760 4980 9824
rect 5044 9760 5060 9824
rect 5124 9760 5140 9824
rect 5204 9760 5210 9824
rect 4894 9759 5210 9760
rect 8842 9824 9158 9825
rect 8842 9760 8848 9824
rect 8912 9760 8928 9824
rect 8992 9760 9008 9824
rect 9072 9760 9088 9824
rect 9152 9760 9158 9824
rect 8842 9759 9158 9760
rect 12790 9824 13106 9825
rect 12790 9760 12796 9824
rect 12860 9760 12876 9824
rect 12940 9760 12956 9824
rect 13020 9760 13036 9824
rect 13100 9760 13106 9824
rect 12790 9759 13106 9760
rect 4061 9754 4127 9757
rect 0 9752 4127 9754
rect 0 9696 4066 9752
rect 4122 9696 4127 9752
rect 0 9694 4127 9696
rect 0 9664 400 9694
rect 4061 9691 4127 9694
rect 6821 9754 6887 9757
rect 7598 9754 7604 9756
rect 6821 9752 7604 9754
rect 6821 9696 6826 9752
rect 6882 9696 7604 9752
rect 6821 9694 7604 9696
rect 6821 9691 6887 9694
rect 7598 9692 7604 9694
rect 7668 9754 7674 9756
rect 7925 9754 7991 9757
rect 9581 9756 9647 9757
rect 9581 9754 9628 9756
rect 7668 9752 7991 9754
rect 7668 9696 7930 9752
rect 7986 9696 7991 9752
rect 7668 9694 7991 9696
rect 9536 9752 9628 9754
rect 9536 9696 9586 9752
rect 9536 9694 9628 9696
rect 7668 9692 7674 9694
rect 7925 9691 7991 9694
rect 9581 9692 9628 9694
rect 9692 9692 9698 9756
rect 10174 9692 10180 9756
rect 10244 9754 10250 9756
rect 11973 9754 12039 9757
rect 10244 9752 12039 9754
rect 10244 9696 11978 9752
rect 12034 9696 12039 9752
rect 10244 9694 12039 9696
rect 10244 9692 10250 9694
rect 9581 9691 9647 9692
rect 11973 9691 12039 9694
rect 15653 9752 15719 9757
rect 15653 9696 15658 9752
rect 15714 9696 15719 9752
rect 15653 9691 15719 9696
rect 4337 9618 4403 9621
rect 11278 9618 11284 9620
rect 4337 9616 11284 9618
rect 4337 9560 4342 9616
rect 4398 9560 11284 9616
rect 4337 9558 11284 9560
rect 4337 9555 4403 9558
rect 11278 9556 11284 9558
rect 11348 9556 11354 9620
rect 11646 9556 11652 9620
rect 11716 9618 11722 9620
rect 11789 9618 11855 9621
rect 11716 9616 11855 9618
rect 11716 9560 11794 9616
rect 11850 9560 11855 9616
rect 11716 9558 11855 9560
rect 11716 9556 11722 9558
rect 11789 9555 11855 9558
rect 11973 9618 12039 9621
rect 15656 9618 15716 9691
rect 11973 9616 15716 9618
rect 11973 9560 11978 9616
rect 12034 9560 15716 9616
rect 11973 9558 15716 9560
rect 11973 9555 12039 9558
rect 2129 9482 2195 9485
rect 3734 9482 3740 9484
rect 2129 9480 3740 9482
rect 2129 9424 2134 9480
rect 2190 9424 3740 9480
rect 2129 9422 3740 9424
rect 2129 9419 2195 9422
rect 3734 9420 3740 9422
rect 3804 9482 3810 9484
rect 10542 9482 10548 9484
rect 3804 9422 10548 9482
rect 3804 9420 3810 9422
rect 10542 9420 10548 9422
rect 10612 9420 10618 9484
rect 10685 9482 10751 9485
rect 13302 9482 13308 9484
rect 10685 9480 13308 9482
rect 10685 9424 10690 9480
rect 10746 9424 13308 9480
rect 10685 9422 13308 9424
rect 10685 9419 10751 9422
rect 13302 9420 13308 9422
rect 13372 9420 13378 9484
rect 13629 9482 13695 9485
rect 16389 9482 16455 9485
rect 13629 9480 16455 9482
rect 13629 9424 13634 9480
rect 13690 9424 16394 9480
rect 16450 9424 16455 9480
rect 13629 9422 16455 9424
rect 13629 9419 13695 9422
rect 16389 9419 16455 9422
rect 6085 9346 6151 9349
rect 6678 9346 6684 9348
rect 6085 9344 6684 9346
rect 6085 9288 6090 9344
rect 6146 9288 6684 9344
rect 6085 9286 6684 9288
rect 6085 9283 6151 9286
rect 6678 9284 6684 9286
rect 6748 9284 6754 9348
rect 12341 9346 12407 9349
rect 14549 9346 14615 9349
rect 12341 9344 14615 9346
rect 12341 9288 12346 9344
rect 12402 9288 14554 9344
rect 14610 9288 14615 9344
rect 12341 9286 14615 9288
rect 12341 9283 12407 9286
rect 14549 9283 14615 9286
rect 2920 9280 3236 9281
rect 2920 9216 2926 9280
rect 2990 9216 3006 9280
rect 3070 9216 3086 9280
rect 3150 9216 3166 9280
rect 3230 9216 3236 9280
rect 2920 9215 3236 9216
rect 6868 9280 7184 9281
rect 6868 9216 6874 9280
rect 6938 9216 6954 9280
rect 7018 9216 7034 9280
rect 7098 9216 7114 9280
rect 7178 9216 7184 9280
rect 6868 9215 7184 9216
rect 10816 9280 11132 9281
rect 10816 9216 10822 9280
rect 10886 9216 10902 9280
rect 10966 9216 10982 9280
rect 11046 9216 11062 9280
rect 11126 9216 11132 9280
rect 10816 9215 11132 9216
rect 14764 9280 15080 9281
rect 14764 9216 14770 9280
rect 14834 9216 14850 9280
rect 14914 9216 14930 9280
rect 14994 9216 15010 9280
rect 15074 9216 15080 9280
rect 14764 9215 15080 9216
rect 9581 9210 9647 9213
rect 7284 9208 9647 9210
rect 7284 9152 9586 9208
rect 9642 9152 9647 9208
rect 7284 9150 9647 9152
rect 6177 9074 6243 9077
rect 7284 9074 7344 9150
rect 9581 9147 9647 9150
rect 11329 9210 11395 9213
rect 14181 9210 14247 9213
rect 11329 9208 14247 9210
rect 11329 9152 11334 9208
rect 11390 9152 14186 9208
rect 14242 9152 14247 9208
rect 11329 9150 14247 9152
rect 11329 9147 11395 9150
rect 14181 9147 14247 9150
rect 6177 9072 7344 9074
rect 6177 9016 6182 9072
rect 6238 9016 7344 9072
rect 6177 9014 7344 9016
rect 8753 9074 8819 9077
rect 13261 9074 13327 9077
rect 13997 9076 14063 9077
rect 13997 9074 14044 9076
rect 8753 9072 13327 9074
rect 8753 9016 8758 9072
rect 8814 9016 13266 9072
rect 13322 9016 13327 9072
rect 8753 9014 13327 9016
rect 13952 9072 14044 9074
rect 13952 9016 14002 9072
rect 13952 9014 14044 9016
rect 6177 9011 6243 9014
rect 8753 9011 8819 9014
rect 13261 9011 13327 9014
rect 13997 9012 14044 9014
rect 14108 9012 14114 9076
rect 14549 9074 14615 9077
rect 15694 9074 15700 9076
rect 14549 9072 15700 9074
rect 14549 9016 14554 9072
rect 14610 9016 15700 9072
rect 14549 9014 15700 9016
rect 13997 9011 14063 9012
rect 14549 9011 14615 9014
rect 15694 9012 15700 9014
rect 15764 9012 15770 9076
rect 6269 8938 6335 8941
rect 12525 8938 12591 8941
rect 6269 8936 12591 8938
rect 6269 8880 6274 8936
rect 6330 8880 12530 8936
rect 12586 8880 12591 8936
rect 6269 8878 12591 8880
rect 6269 8875 6335 8878
rect 12525 8875 12591 8878
rect 12985 8938 13051 8941
rect 12985 8936 13554 8938
rect 12985 8880 12990 8936
rect 13046 8880 13554 8936
rect 12985 8878 13554 8880
rect 12985 8875 13051 8878
rect 6729 8802 6795 8805
rect 8661 8802 8727 8805
rect 6729 8800 8727 8802
rect 6729 8744 6734 8800
rect 6790 8744 8666 8800
rect 8722 8744 8727 8800
rect 6729 8742 8727 8744
rect 6729 8739 6795 8742
rect 8661 8739 8727 8742
rect 10542 8740 10548 8804
rect 10612 8802 10618 8804
rect 13494 8802 13554 8878
rect 13854 8876 13860 8940
rect 13924 8938 13930 8940
rect 15101 8938 15167 8941
rect 15377 8938 15443 8941
rect 13924 8936 15167 8938
rect 13924 8880 15106 8936
rect 15162 8880 15167 8936
rect 13924 8878 15167 8880
rect 13924 8876 13930 8878
rect 15101 8875 15167 8878
rect 15334 8936 15443 8938
rect 15334 8880 15382 8936
rect 15438 8880 15443 8936
rect 15334 8875 15443 8880
rect 14733 8802 14799 8805
rect 10612 8742 12404 8802
rect 13494 8800 14799 8802
rect 13494 8744 14738 8800
rect 14794 8744 14799 8800
rect 13494 8742 14799 8744
rect 10612 8740 10618 8742
rect 4894 8736 5210 8737
rect 4894 8672 4900 8736
rect 4964 8672 4980 8736
rect 5044 8672 5060 8736
rect 5124 8672 5140 8736
rect 5204 8672 5210 8736
rect 4894 8671 5210 8672
rect 8842 8736 9158 8737
rect 8842 8672 8848 8736
rect 8912 8672 8928 8736
rect 8992 8672 9008 8736
rect 9072 8672 9088 8736
rect 9152 8672 9158 8736
rect 8842 8671 9158 8672
rect 2681 8666 2747 8669
rect 4429 8666 4495 8669
rect 2681 8664 4495 8666
rect 2681 8608 2686 8664
rect 2742 8608 4434 8664
rect 4490 8608 4495 8664
rect 2681 8606 4495 8608
rect 2681 8603 2747 8606
rect 4429 8603 4495 8606
rect 5441 8666 5507 8669
rect 8661 8666 8727 8669
rect 5441 8664 8727 8666
rect 5441 8608 5446 8664
rect 5502 8608 8666 8664
rect 8722 8608 8727 8664
rect 5441 8606 8727 8608
rect 5441 8603 5507 8606
rect 8661 8603 8727 8606
rect 9581 8666 9647 8669
rect 10869 8666 10935 8669
rect 9581 8664 10935 8666
rect 9581 8608 9586 8664
rect 9642 8608 10874 8664
rect 10930 8608 10935 8664
rect 9581 8606 10935 8608
rect 9581 8603 9647 8606
rect 10869 8603 10935 8606
rect 3601 8530 3667 8533
rect 4061 8530 4127 8533
rect 3601 8528 4127 8530
rect 3601 8472 3606 8528
rect 3662 8472 4066 8528
rect 4122 8472 4127 8528
rect 3601 8470 4127 8472
rect 3601 8467 3667 8470
rect 4061 8467 4127 8470
rect 4337 8530 4403 8533
rect 12344 8530 12404 8742
rect 14733 8739 14799 8742
rect 12790 8736 13106 8737
rect 12790 8672 12796 8736
rect 12860 8672 12876 8736
rect 12940 8672 12956 8736
rect 13020 8672 13036 8736
rect 13100 8672 13106 8736
rect 12790 8671 13106 8672
rect 12525 8668 12591 8669
rect 12525 8664 12572 8668
rect 12636 8666 12642 8668
rect 12525 8608 12530 8664
rect 12525 8604 12572 8608
rect 12636 8606 12682 8666
rect 12636 8604 12642 8606
rect 13302 8604 13308 8668
rect 13372 8666 13378 8668
rect 13721 8666 13787 8669
rect 14406 8666 14412 8668
rect 13372 8664 13787 8666
rect 13372 8608 13726 8664
rect 13782 8608 13787 8664
rect 13372 8606 13787 8608
rect 13372 8604 13378 8606
rect 12525 8603 12591 8604
rect 13721 8603 13787 8606
rect 13862 8606 14412 8666
rect 13721 8530 13787 8533
rect 13862 8530 13922 8606
rect 14406 8604 14412 8606
rect 14476 8604 14482 8668
rect 15334 8666 15394 8875
rect 15150 8606 15394 8666
rect 4337 8528 12266 8530
rect 4337 8472 4342 8528
rect 4398 8472 12266 8528
rect 4337 8470 12266 8472
rect 12344 8528 13922 8530
rect 12344 8472 13726 8528
rect 13782 8472 13922 8528
rect 12344 8470 13922 8472
rect 4337 8467 4403 8470
rect 4061 8394 4127 8397
rect 4470 8394 4476 8396
rect 4061 8392 4476 8394
rect 4061 8336 4066 8392
rect 4122 8336 4476 8392
rect 4061 8334 4476 8336
rect 4061 8331 4127 8334
rect 4470 8332 4476 8334
rect 4540 8332 4546 8396
rect 4654 8332 4660 8396
rect 4724 8394 4730 8396
rect 5073 8394 5139 8397
rect 4724 8392 5139 8394
rect 4724 8336 5078 8392
rect 5134 8336 5139 8392
rect 4724 8334 5139 8336
rect 4724 8332 4730 8334
rect 5073 8331 5139 8334
rect 8293 8394 8359 8397
rect 12206 8396 12266 8470
rect 13721 8467 13787 8470
rect 14406 8468 14412 8532
rect 14476 8530 14482 8532
rect 14733 8530 14799 8533
rect 15150 8530 15210 8606
rect 16062 8530 16068 8532
rect 14476 8528 15210 8530
rect 14476 8472 14738 8528
rect 14794 8472 15210 8528
rect 14476 8470 15210 8472
rect 15288 8470 16068 8530
rect 14476 8468 14482 8470
rect 14733 8467 14799 8470
rect 11646 8394 11652 8396
rect 8293 8392 11652 8394
rect 8293 8336 8298 8392
rect 8354 8336 11652 8392
rect 8293 8334 11652 8336
rect 8293 8331 8359 8334
rect 11646 8332 11652 8334
rect 11716 8332 11722 8396
rect 12198 8332 12204 8396
rect 12268 8394 12274 8396
rect 14825 8394 14891 8397
rect 12268 8392 14891 8394
rect 12268 8336 14830 8392
rect 14886 8336 14891 8392
rect 12268 8334 14891 8336
rect 12268 8332 12274 8334
rect 14825 8331 14891 8334
rect 15101 8394 15167 8397
rect 15288 8394 15348 8470
rect 16062 8468 16068 8470
rect 16132 8468 16138 8532
rect 15745 8396 15811 8397
rect 15101 8392 15348 8394
rect 15101 8336 15106 8392
rect 15162 8336 15348 8392
rect 15101 8334 15348 8336
rect 15101 8331 15167 8334
rect 15694 8332 15700 8396
rect 15764 8394 15811 8396
rect 15764 8392 15856 8394
rect 15806 8336 15856 8392
rect 15764 8334 15856 8336
rect 15764 8332 15811 8334
rect 15745 8331 15811 8332
rect 0 8258 400 8288
rect 473 8258 539 8261
rect 0 8256 539 8258
rect 0 8200 478 8256
rect 534 8200 539 8256
rect 0 8198 539 8200
rect 0 8168 400 8198
rect 473 8195 539 8198
rect 8150 8196 8156 8260
rect 8220 8258 8226 8260
rect 8753 8258 8819 8261
rect 8220 8256 8819 8258
rect 8220 8200 8758 8256
rect 8814 8200 8819 8256
rect 8220 8198 8819 8200
rect 8220 8196 8226 8198
rect 8753 8195 8819 8198
rect 9029 8258 9095 8261
rect 9305 8258 9371 8261
rect 9622 8258 9628 8260
rect 9029 8256 9628 8258
rect 9029 8200 9034 8256
rect 9090 8200 9310 8256
rect 9366 8200 9628 8256
rect 9029 8198 9628 8200
rect 9029 8195 9095 8198
rect 9305 8195 9371 8198
rect 9622 8196 9628 8198
rect 9692 8196 9698 8260
rect 11237 8258 11303 8261
rect 14222 8258 14228 8260
rect 11237 8256 14228 8258
rect 11237 8200 11242 8256
rect 11298 8200 14228 8256
rect 11237 8198 14228 8200
rect 11237 8195 11303 8198
rect 14222 8196 14228 8198
rect 14292 8196 14298 8260
rect 2920 8192 3236 8193
rect 2920 8128 2926 8192
rect 2990 8128 3006 8192
rect 3070 8128 3086 8192
rect 3150 8128 3166 8192
rect 3230 8128 3236 8192
rect 2920 8127 3236 8128
rect 6868 8192 7184 8193
rect 6868 8128 6874 8192
rect 6938 8128 6954 8192
rect 7018 8128 7034 8192
rect 7098 8128 7114 8192
rect 7178 8128 7184 8192
rect 6868 8127 7184 8128
rect 10816 8192 11132 8193
rect 10816 8128 10822 8192
rect 10886 8128 10902 8192
rect 10966 8128 10982 8192
rect 11046 8128 11062 8192
rect 11126 8128 11132 8192
rect 10816 8127 11132 8128
rect 14764 8192 15080 8193
rect 14764 8128 14770 8192
rect 14834 8128 14850 8192
rect 14914 8128 14930 8192
rect 14994 8128 15010 8192
rect 15074 8128 15080 8192
rect 14764 8127 15080 8128
rect 7598 8060 7604 8124
rect 7668 8122 7674 8124
rect 9806 8122 9812 8124
rect 7668 8062 9812 8122
rect 7668 8060 7674 8062
rect 9806 8060 9812 8062
rect 9876 8122 9882 8124
rect 9876 8062 10610 8122
rect 9876 8060 9882 8062
rect 5758 7924 5764 7988
rect 5828 7986 5834 7988
rect 6177 7986 6243 7989
rect 5828 7984 6243 7986
rect 5828 7928 6182 7984
rect 6238 7928 6243 7984
rect 5828 7926 6243 7928
rect 5828 7924 5834 7926
rect 6177 7923 6243 7926
rect 6545 7986 6611 7989
rect 9213 7986 9279 7989
rect 6545 7984 9279 7986
rect 6545 7928 6550 7984
rect 6606 7928 9218 7984
rect 9274 7928 9279 7984
rect 6545 7926 9279 7928
rect 6545 7923 6611 7926
rect 9213 7923 9279 7926
rect 9622 7924 9628 7988
rect 9692 7986 9698 7988
rect 10550 7986 10610 8062
rect 11830 8060 11836 8124
rect 11900 8122 11906 8124
rect 12382 8122 12388 8124
rect 11900 8062 12388 8122
rect 11900 8060 11906 8062
rect 12382 8060 12388 8062
rect 12452 8060 12458 8124
rect 13905 8122 13971 8125
rect 14089 8122 14155 8125
rect 13905 8120 14155 8122
rect 13905 8064 13910 8120
rect 13966 8064 14094 8120
rect 14150 8064 14155 8120
rect 13905 8062 14155 8064
rect 13905 8059 13971 8062
rect 14089 8059 14155 8062
rect 10777 7986 10843 7989
rect 9692 7926 10058 7986
rect 10550 7984 10843 7986
rect 10550 7928 10782 7984
rect 10838 7928 10843 7984
rect 10550 7926 10843 7928
rect 9692 7924 9698 7926
rect 4286 7788 4292 7852
rect 4356 7850 4362 7852
rect 4797 7850 4863 7853
rect 4356 7848 9322 7850
rect 4356 7792 4802 7848
rect 4858 7792 9322 7848
rect 4356 7790 9322 7792
rect 4356 7788 4362 7790
rect 4797 7787 4863 7790
rect 5574 7652 5580 7716
rect 5644 7714 5650 7716
rect 8569 7714 8635 7717
rect 5644 7712 8635 7714
rect 5644 7656 8574 7712
rect 8630 7656 8635 7712
rect 5644 7654 8635 7656
rect 5644 7652 5650 7654
rect 8569 7651 8635 7654
rect 4894 7648 5210 7649
rect 4894 7584 4900 7648
rect 4964 7584 4980 7648
rect 5044 7584 5060 7648
rect 5124 7584 5140 7648
rect 5204 7584 5210 7648
rect 4894 7583 5210 7584
rect 8842 7648 9158 7649
rect 8842 7584 8848 7648
rect 8912 7584 8928 7648
rect 8992 7584 9008 7648
rect 9072 7584 9088 7648
rect 9152 7584 9158 7648
rect 8842 7583 9158 7584
rect 6177 7578 6243 7581
rect 9262 7578 9322 7790
rect 9622 7788 9628 7852
rect 9692 7850 9698 7852
rect 9857 7850 9923 7853
rect 9692 7848 9923 7850
rect 9692 7792 9862 7848
rect 9918 7792 9923 7848
rect 9692 7790 9923 7792
rect 9998 7850 10058 7926
rect 10777 7923 10843 7926
rect 12382 7924 12388 7988
rect 12452 7986 12458 7988
rect 12709 7986 12775 7989
rect 12452 7984 12775 7986
rect 12452 7928 12714 7984
rect 12770 7928 12775 7984
rect 12452 7926 12775 7928
rect 12452 7924 12458 7926
rect 12709 7923 12775 7926
rect 12893 7986 12959 7989
rect 15101 7986 15167 7989
rect 12893 7984 15167 7986
rect 12893 7928 12898 7984
rect 12954 7928 15106 7984
rect 15162 7928 15167 7984
rect 12893 7926 15167 7928
rect 12893 7923 12959 7926
rect 15101 7923 15167 7926
rect 10961 7850 11027 7853
rect 11421 7852 11487 7853
rect 11421 7850 11468 7852
rect 9998 7848 11027 7850
rect 9998 7792 10966 7848
rect 11022 7792 11027 7848
rect 9998 7790 11027 7792
rect 11376 7848 11468 7850
rect 11376 7792 11426 7848
rect 11376 7790 11468 7792
rect 9692 7788 9698 7790
rect 9857 7787 9923 7790
rect 10961 7787 11027 7790
rect 11421 7788 11468 7790
rect 11532 7788 11538 7852
rect 11881 7850 11947 7853
rect 12198 7850 12204 7852
rect 11881 7848 12204 7850
rect 11881 7792 11886 7848
rect 11942 7792 12204 7848
rect 11881 7790 12204 7792
rect 11421 7787 11487 7788
rect 11881 7787 11947 7790
rect 12198 7788 12204 7790
rect 12268 7788 12274 7852
rect 12433 7850 12499 7853
rect 13813 7852 13879 7853
rect 12566 7850 12572 7852
rect 12433 7848 12572 7850
rect 12433 7792 12438 7848
rect 12494 7792 12572 7848
rect 12433 7790 12572 7792
rect 12433 7787 12499 7790
rect 12566 7788 12572 7790
rect 12636 7788 12642 7852
rect 13813 7848 13860 7852
rect 13924 7850 13930 7852
rect 13813 7792 13818 7848
rect 13813 7788 13860 7792
rect 13924 7790 13970 7850
rect 14641 7848 14707 7853
rect 14641 7792 14646 7848
rect 14702 7792 14707 7848
rect 13924 7788 13930 7790
rect 13813 7787 13879 7788
rect 14641 7787 14707 7792
rect 9438 7652 9444 7716
rect 9508 7714 9514 7716
rect 12433 7714 12499 7717
rect 14644 7714 14704 7787
rect 9508 7712 12499 7714
rect 9508 7656 12438 7712
rect 12494 7656 12499 7712
rect 9508 7654 12499 7656
rect 9508 7652 9514 7654
rect 12433 7651 12499 7654
rect 13172 7654 14704 7714
rect 12790 7648 13106 7649
rect 12790 7584 12796 7648
rect 12860 7584 12876 7648
rect 12940 7584 12956 7648
rect 13020 7584 13036 7648
rect 13100 7584 13106 7648
rect 12790 7583 13106 7584
rect 6177 7576 8172 7578
rect 6177 7520 6182 7576
rect 6238 7520 8172 7576
rect 6177 7518 8172 7520
rect 9262 7518 12634 7578
rect 6177 7515 6243 7518
rect 4102 7380 4108 7444
rect 4172 7442 4178 7444
rect 5625 7442 5691 7445
rect 4172 7440 5691 7442
rect 4172 7384 5630 7440
rect 5686 7384 5691 7440
rect 4172 7382 5691 7384
rect 4172 7380 4178 7382
rect 5625 7379 5691 7382
rect 7005 7442 7071 7445
rect 7925 7442 7991 7445
rect 7005 7440 7991 7442
rect 7005 7384 7010 7440
rect 7066 7384 7930 7440
rect 7986 7384 7991 7440
rect 7005 7382 7991 7384
rect 8112 7442 8172 7518
rect 9857 7442 9923 7445
rect 9990 7442 9996 7444
rect 8112 7440 9996 7442
rect 8112 7384 9862 7440
rect 9918 7384 9996 7440
rect 8112 7382 9996 7384
rect 7005 7379 7071 7382
rect 7925 7379 7991 7382
rect 9857 7379 9923 7382
rect 9990 7380 9996 7382
rect 10060 7380 10066 7444
rect 10961 7442 11027 7445
rect 12574 7442 12634 7518
rect 13172 7442 13232 7654
rect 13905 7578 13971 7581
rect 16614 7578 16620 7580
rect 13905 7576 16620 7578
rect 13905 7520 13910 7576
rect 13966 7520 16620 7576
rect 13905 7518 16620 7520
rect 13905 7515 13971 7518
rect 16614 7516 16620 7518
rect 16684 7516 16690 7580
rect 10961 7440 11852 7442
rect 10961 7384 10966 7440
rect 11022 7384 11852 7440
rect 10961 7382 11852 7384
rect 12574 7382 13232 7442
rect 16297 7440 16363 7445
rect 16297 7384 16302 7440
rect 16358 7384 16363 7440
rect 10961 7379 11027 7382
rect 3601 7306 3667 7309
rect 11605 7306 11671 7309
rect 3601 7304 11671 7306
rect 3601 7248 3606 7304
rect 3662 7248 11610 7304
rect 11666 7248 11671 7304
rect 3601 7246 11671 7248
rect 11792 7306 11852 7382
rect 16297 7379 16363 7384
rect 13905 7306 13971 7309
rect 11792 7304 13971 7306
rect 11792 7248 13910 7304
rect 13966 7248 13971 7304
rect 11792 7246 13971 7248
rect 3601 7243 3667 7246
rect 11605 7243 11671 7246
rect 13905 7243 13971 7246
rect 8017 7170 8083 7173
rect 9121 7170 9187 7173
rect 8017 7168 9187 7170
rect 8017 7112 8022 7168
rect 8078 7112 9126 7168
rect 9182 7112 9187 7168
rect 8017 7110 9187 7112
rect 8017 7107 8083 7110
rect 9121 7107 9187 7110
rect 9765 7172 9831 7173
rect 9765 7168 9812 7172
rect 9876 7170 9882 7172
rect 9765 7112 9770 7168
rect 9765 7108 9812 7112
rect 9876 7110 9922 7170
rect 9876 7108 9882 7110
rect 11278 7108 11284 7172
rect 11348 7170 11354 7172
rect 12433 7170 12499 7173
rect 11348 7168 12499 7170
rect 11348 7112 12438 7168
rect 12494 7112 12499 7168
rect 11348 7110 12499 7112
rect 11348 7108 11354 7110
rect 9765 7107 9831 7108
rect 12433 7107 12499 7110
rect 2920 7104 3236 7105
rect 2920 7040 2926 7104
rect 2990 7040 3006 7104
rect 3070 7040 3086 7104
rect 3150 7040 3166 7104
rect 3230 7040 3236 7104
rect 2920 7039 3236 7040
rect 6868 7104 7184 7105
rect 6868 7040 6874 7104
rect 6938 7040 6954 7104
rect 7018 7040 7034 7104
rect 7098 7040 7114 7104
rect 7178 7040 7184 7104
rect 6868 7039 7184 7040
rect 10816 7104 11132 7105
rect 10816 7040 10822 7104
rect 10886 7040 10902 7104
rect 10966 7040 10982 7104
rect 11046 7040 11062 7104
rect 11126 7040 11132 7104
rect 10816 7039 11132 7040
rect 14764 7104 15080 7105
rect 14764 7040 14770 7104
rect 14834 7040 14850 7104
rect 14914 7040 14930 7104
rect 14994 7040 15010 7104
rect 15074 7040 15080 7104
rect 14764 7039 15080 7040
rect 8661 7034 8727 7037
rect 9254 7034 9260 7036
rect 8661 7032 9260 7034
rect 8661 6976 8666 7032
rect 8722 6976 9260 7032
rect 8661 6974 9260 6976
rect 8661 6971 8727 6974
rect 9254 6972 9260 6974
rect 9324 6972 9330 7036
rect 9765 7034 9831 7037
rect 10041 7034 10107 7037
rect 9765 7032 10107 7034
rect 9765 6976 9770 7032
rect 9826 6976 10046 7032
rect 10102 6976 10107 7032
rect 9765 6974 10107 6976
rect 9765 6971 9831 6974
rect 10041 6971 10107 6974
rect 11237 7034 11303 7037
rect 11237 7032 13692 7034
rect 11237 6976 11242 7032
rect 11298 6976 13692 7032
rect 11237 6974 13692 6976
rect 11237 6971 11303 6974
rect 2681 6900 2747 6901
rect 2630 6898 2636 6900
rect 2590 6838 2636 6898
rect 2700 6896 2747 6900
rect 2742 6840 2747 6896
rect 2630 6836 2636 6838
rect 2700 6836 2747 6840
rect 2681 6835 2747 6836
rect 3509 6898 3575 6901
rect 11053 6898 11119 6901
rect 3509 6896 11119 6898
rect 3509 6840 3514 6896
rect 3570 6840 11058 6896
rect 11114 6840 11119 6896
rect 3509 6838 11119 6840
rect 3509 6835 3575 6838
rect 11053 6835 11119 6838
rect 11278 6836 11284 6900
rect 11348 6898 11354 6900
rect 13445 6898 13511 6901
rect 11348 6896 13511 6898
rect 11348 6840 13450 6896
rect 13506 6840 13511 6896
rect 11348 6838 13511 6840
rect 13632 6898 13692 6974
rect 16300 6901 16360 7379
rect 15326 6898 15332 6900
rect 13632 6838 15332 6898
rect 11348 6836 11354 6838
rect 13445 6835 13511 6838
rect 15326 6836 15332 6838
rect 15396 6898 15402 6900
rect 15561 6898 15627 6901
rect 15396 6896 15627 6898
rect 15396 6840 15566 6896
rect 15622 6840 15627 6896
rect 15396 6838 15627 6840
rect 15396 6836 15402 6838
rect 15561 6835 15627 6838
rect 16297 6896 16363 6901
rect 16297 6840 16302 6896
rect 16358 6840 16363 6896
rect 16297 6835 16363 6840
rect 0 6762 400 6792
rect 8109 6762 8175 6765
rect 9949 6762 10015 6765
rect 0 6760 8175 6762
rect 0 6704 8114 6760
rect 8170 6704 8175 6760
rect 0 6702 8175 6704
rect 0 6672 400 6702
rect 8109 6699 8175 6702
rect 8250 6760 10015 6762
rect 8250 6704 9954 6760
rect 10010 6704 10015 6760
rect 8250 6702 10015 6704
rect 6269 6626 6335 6629
rect 8250 6626 8310 6702
rect 9949 6699 10015 6702
rect 10174 6700 10180 6764
rect 10244 6762 10250 6764
rect 17677 6762 17743 6765
rect 10244 6760 17743 6762
rect 10244 6704 17682 6760
rect 17738 6704 17743 6760
rect 10244 6702 17743 6704
rect 10244 6700 10250 6702
rect 17677 6699 17743 6702
rect 6269 6624 8310 6626
rect 6269 6568 6274 6624
rect 6330 6568 8310 6624
rect 6269 6566 8310 6568
rect 9581 6626 9647 6629
rect 10869 6626 10935 6629
rect 9581 6624 10935 6626
rect 9581 6568 9586 6624
rect 9642 6568 10874 6624
rect 10930 6568 10935 6624
rect 9581 6566 10935 6568
rect 6269 6563 6335 6566
rect 9581 6563 9647 6566
rect 10869 6563 10935 6566
rect 11053 6626 11119 6629
rect 12617 6626 12683 6629
rect 11053 6624 12683 6626
rect 11053 6568 11058 6624
rect 11114 6568 12622 6624
rect 12678 6568 12683 6624
rect 11053 6566 12683 6568
rect 11053 6563 11119 6566
rect 12617 6563 12683 6566
rect 13261 6626 13327 6629
rect 15326 6626 15332 6628
rect 13261 6624 15332 6626
rect 13261 6568 13266 6624
rect 13322 6568 15332 6624
rect 13261 6566 15332 6568
rect 13261 6563 13327 6566
rect 15326 6564 15332 6566
rect 15396 6626 15402 6628
rect 15694 6626 15700 6628
rect 15396 6566 15700 6626
rect 15396 6564 15402 6566
rect 15694 6564 15700 6566
rect 15764 6564 15770 6628
rect 4894 6560 5210 6561
rect 4894 6496 4900 6560
rect 4964 6496 4980 6560
rect 5044 6496 5060 6560
rect 5124 6496 5140 6560
rect 5204 6496 5210 6560
rect 4894 6495 5210 6496
rect 8842 6560 9158 6561
rect 8842 6496 8848 6560
rect 8912 6496 8928 6560
rect 8992 6496 9008 6560
rect 9072 6496 9088 6560
rect 9152 6496 9158 6560
rect 8842 6495 9158 6496
rect 12790 6560 13106 6561
rect 12790 6496 12796 6560
rect 12860 6496 12876 6560
rect 12940 6496 12956 6560
rect 13020 6496 13036 6560
rect 13100 6496 13106 6560
rect 12790 6495 13106 6496
rect 7189 6490 7255 6493
rect 7557 6490 7623 6493
rect 8201 6492 8267 6493
rect 8150 6490 8156 6492
rect 7189 6488 7623 6490
rect 7189 6432 7194 6488
rect 7250 6432 7562 6488
rect 7618 6432 7623 6488
rect 7189 6430 7623 6432
rect 8110 6430 8156 6490
rect 8220 6488 8267 6492
rect 8262 6432 8267 6488
rect 7189 6427 7255 6430
rect 7557 6427 7623 6430
rect 8150 6428 8156 6430
rect 8220 6428 8267 6432
rect 8201 6427 8267 6428
rect 9949 6490 10015 6493
rect 11973 6490 12039 6493
rect 9949 6488 12039 6490
rect 9949 6432 9954 6488
rect 10010 6432 11978 6488
rect 12034 6432 12039 6488
rect 9949 6430 12039 6432
rect 9949 6427 10015 6430
rect 11973 6427 12039 6430
rect 13537 6490 13603 6493
rect 13670 6490 13676 6492
rect 13537 6488 13676 6490
rect 13537 6432 13542 6488
rect 13598 6432 13676 6488
rect 13537 6430 13676 6432
rect 13537 6427 13603 6430
rect 13670 6428 13676 6430
rect 13740 6428 13746 6492
rect 3693 6352 3759 6357
rect 3693 6296 3698 6352
rect 3754 6296 3759 6352
rect 3693 6291 3759 6296
rect 7097 6354 7163 6357
rect 8518 6354 8524 6356
rect 7097 6352 8524 6354
rect 7097 6296 7102 6352
rect 7158 6296 8524 6352
rect 7097 6294 8524 6296
rect 7097 6291 7163 6294
rect 8518 6292 8524 6294
rect 8588 6292 8594 6356
rect 8661 6354 8727 6357
rect 11053 6354 11119 6357
rect 8661 6352 11119 6354
rect 8661 6296 8666 6352
rect 8722 6296 11058 6352
rect 11114 6296 11119 6352
rect 8661 6294 11119 6296
rect 8661 6291 8727 6294
rect 2313 6218 2379 6221
rect 3696 6218 3756 6291
rect 9952 6260 10058 6294
rect 11053 6291 11119 6294
rect 11605 6354 11671 6357
rect 12382 6354 12388 6356
rect 11605 6352 12388 6354
rect 11605 6296 11610 6352
rect 11666 6296 12388 6352
rect 11605 6294 12388 6296
rect 11605 6291 11671 6294
rect 12382 6292 12388 6294
rect 12452 6292 12458 6356
rect 12801 6354 12867 6357
rect 13854 6354 13860 6356
rect 12801 6352 13860 6354
rect 12801 6296 12806 6352
rect 12862 6296 13860 6352
rect 12801 6294 13860 6296
rect 12801 6291 12867 6294
rect 13854 6292 13860 6294
rect 13924 6354 13930 6356
rect 15377 6354 15443 6357
rect 13924 6352 15443 6354
rect 13924 6296 15382 6352
rect 15438 6296 15443 6352
rect 13924 6294 15443 6296
rect 13924 6292 13930 6294
rect 15377 6291 15443 6294
rect 2313 6216 3756 6218
rect 2313 6160 2318 6216
rect 2374 6160 3756 6216
rect 2313 6158 3756 6160
rect 2313 6155 2379 6158
rect 3696 6082 3756 6158
rect 4061 6218 4127 6221
rect 9397 6218 9463 6221
rect 4061 6216 9463 6218
rect 4061 6160 4066 6216
rect 4122 6160 9402 6216
rect 9458 6160 9463 6216
rect 4061 6158 9463 6160
rect 4061 6155 4127 6158
rect 9397 6155 9463 6158
rect 10409 6218 10475 6221
rect 16246 6218 16252 6220
rect 10409 6216 16252 6218
rect 10409 6160 10414 6216
rect 10470 6160 16252 6216
rect 10409 6158 16252 6160
rect 10409 6155 10475 6158
rect 16246 6156 16252 6158
rect 16316 6156 16322 6220
rect 5533 6082 5599 6085
rect 3696 6080 5599 6082
rect 3696 6024 5538 6080
rect 5594 6024 5599 6080
rect 3696 6022 5599 6024
rect 5533 6019 5599 6022
rect 7373 6082 7439 6085
rect 10317 6082 10383 6085
rect 7373 6080 10748 6082
rect 7373 6024 7378 6080
rect 7434 6024 10322 6080
rect 10378 6024 10748 6080
rect 7373 6022 10748 6024
rect 7373 6019 7439 6022
rect 10317 6019 10383 6022
rect 2920 6016 3236 6017
rect 2920 5952 2926 6016
rect 2990 5952 3006 6016
rect 3070 5952 3086 6016
rect 3150 5952 3166 6016
rect 3230 5952 3236 6016
rect 2920 5951 3236 5952
rect 6868 6016 7184 6017
rect 6868 5952 6874 6016
rect 6938 5952 6954 6016
rect 7018 5952 7034 6016
rect 7098 5952 7114 6016
rect 7178 5952 7184 6016
rect 6868 5951 7184 5952
rect 8845 5946 8911 5949
rect 9213 5946 9279 5949
rect 9622 5946 9628 5948
rect 8845 5944 9138 5946
rect 8845 5888 8850 5944
rect 8906 5888 9138 5944
rect 8845 5886 9138 5888
rect 8845 5883 8911 5886
rect 2681 5810 2747 5813
rect 2681 5808 5550 5810
rect 2681 5752 2686 5808
rect 2742 5752 5550 5808
rect 2681 5750 5550 5752
rect 2681 5747 2747 5750
rect 4061 5676 4127 5677
rect 4061 5674 4108 5676
rect 4016 5672 4108 5674
rect 4016 5616 4066 5672
rect 4016 5614 4108 5616
rect 4061 5612 4108 5614
rect 4172 5612 4178 5676
rect 5490 5674 5550 5750
rect 6310 5748 6316 5812
rect 6380 5810 6386 5812
rect 8937 5810 9003 5813
rect 6380 5808 9003 5810
rect 6380 5752 8942 5808
rect 8998 5752 9003 5808
rect 6380 5750 9003 5752
rect 9078 5810 9138 5886
rect 9213 5944 9628 5946
rect 9213 5888 9218 5944
rect 9274 5888 9628 5944
rect 9213 5886 9628 5888
rect 9213 5883 9279 5886
rect 9622 5884 9628 5886
rect 9692 5884 9698 5948
rect 9765 5946 9831 5949
rect 10501 5946 10567 5949
rect 9765 5944 10567 5946
rect 9765 5888 9770 5944
rect 9826 5888 10506 5944
rect 10562 5888 10567 5944
rect 9765 5886 10567 5888
rect 9765 5883 9831 5886
rect 10501 5883 10567 5886
rect 10688 5844 10748 6022
rect 11462 6020 11468 6084
rect 11532 6082 11538 6084
rect 14181 6082 14247 6085
rect 11532 6080 14247 6082
rect 11532 6024 14186 6080
rect 14242 6024 14247 6080
rect 11532 6022 14247 6024
rect 11532 6020 11538 6022
rect 14181 6019 14247 6022
rect 10816 6016 11132 6017
rect 10816 5952 10822 6016
rect 10886 5952 10902 6016
rect 10966 5952 10982 6016
rect 11046 5952 11062 6016
rect 11126 5952 11132 6016
rect 10816 5951 11132 5952
rect 14764 6016 15080 6017
rect 14764 5952 14770 6016
rect 14834 5952 14850 6016
rect 14914 5952 14930 6016
rect 14994 5952 15010 6016
rect 15074 5952 15080 6016
rect 14764 5951 15080 5952
rect 11605 5946 11671 5949
rect 14406 5946 14412 5948
rect 11605 5944 14412 5946
rect 11605 5888 11610 5944
rect 11666 5888 14412 5944
rect 11605 5886 14412 5888
rect 11605 5883 11671 5886
rect 14406 5884 14412 5886
rect 14476 5884 14482 5948
rect 15193 5944 15259 5949
rect 15193 5888 15198 5944
rect 15254 5888 15259 5944
rect 15193 5883 15259 5888
rect 10225 5810 10291 5813
rect 9078 5808 10291 5810
rect 9078 5752 10230 5808
rect 10286 5752 10291 5808
rect 10688 5810 10794 5844
rect 11053 5810 11119 5813
rect 10688 5808 11119 5810
rect 10688 5784 11058 5808
rect 9078 5750 10291 5752
rect 10734 5752 11058 5784
rect 11114 5752 11119 5808
rect 10734 5750 11119 5752
rect 6380 5748 6386 5750
rect 8937 5747 9003 5750
rect 10225 5747 10291 5750
rect 11053 5747 11119 5750
rect 11881 5810 11947 5813
rect 13169 5810 13235 5813
rect 11881 5808 13235 5810
rect 11881 5752 11886 5808
rect 11942 5752 13174 5808
rect 13230 5752 13235 5808
rect 11881 5750 13235 5752
rect 11881 5747 11947 5750
rect 13169 5747 13235 5750
rect 13353 5810 13419 5813
rect 13670 5810 13676 5812
rect 13353 5808 13676 5810
rect 13353 5752 13358 5808
rect 13414 5752 13676 5808
rect 13353 5750 13676 5752
rect 13353 5747 13419 5750
rect 13670 5748 13676 5750
rect 13740 5748 13746 5812
rect 14457 5810 14523 5813
rect 15196 5810 15256 5883
rect 14457 5808 15256 5810
rect 14457 5752 14462 5808
rect 14518 5752 15256 5808
rect 14457 5750 15256 5752
rect 14457 5747 14523 5750
rect 9305 5674 9371 5677
rect 10501 5674 10567 5677
rect 5490 5672 10567 5674
rect 5490 5616 9310 5672
rect 9366 5616 10506 5672
rect 10562 5616 10567 5672
rect 5490 5614 10567 5616
rect 4061 5611 4127 5612
rect 9305 5611 9371 5614
rect 10501 5611 10567 5614
rect 10777 5674 10843 5677
rect 13356 5674 13416 5747
rect 10777 5672 13416 5674
rect 10777 5616 10782 5672
rect 10838 5616 13416 5672
rect 10777 5614 13416 5616
rect 10777 5611 10843 5614
rect 5533 5538 5599 5541
rect 8293 5538 8359 5541
rect 5533 5536 8359 5538
rect 5533 5480 5538 5536
rect 5594 5480 8298 5536
rect 8354 5480 8359 5536
rect 5533 5478 8359 5480
rect 5533 5475 5599 5478
rect 8293 5475 8359 5478
rect 9622 5476 9628 5540
rect 9692 5538 9698 5540
rect 10358 5538 10364 5540
rect 9692 5478 10364 5538
rect 9692 5476 9698 5478
rect 10358 5476 10364 5478
rect 10428 5476 10434 5540
rect 10593 5538 10659 5541
rect 11462 5538 11468 5540
rect 10593 5536 11468 5538
rect 10593 5480 10598 5536
rect 10654 5480 11468 5536
rect 10593 5478 11468 5480
rect 10593 5475 10659 5478
rect 11462 5476 11468 5478
rect 11532 5476 11538 5540
rect 11881 5538 11947 5541
rect 12198 5538 12204 5540
rect 11700 5536 11947 5538
rect 11700 5480 11886 5536
rect 11942 5480 11947 5536
rect 11700 5478 11947 5480
rect 4894 5472 5210 5473
rect 4894 5408 4900 5472
rect 4964 5408 4980 5472
rect 5044 5408 5060 5472
rect 5124 5408 5140 5472
rect 5204 5408 5210 5472
rect 4894 5407 5210 5408
rect 8842 5472 9158 5473
rect 8842 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9008 5472
rect 9072 5408 9088 5472
rect 9152 5408 9158 5472
rect 8842 5407 9158 5408
rect 6453 5402 6519 5405
rect 6729 5402 6795 5405
rect 6453 5400 6795 5402
rect 6453 5344 6458 5400
rect 6514 5344 6734 5400
rect 6790 5344 6795 5400
rect 6453 5342 6795 5344
rect 6453 5339 6519 5342
rect 6729 5339 6795 5342
rect 7005 5402 7071 5405
rect 7966 5402 7972 5404
rect 7005 5400 7972 5402
rect 7005 5344 7010 5400
rect 7066 5344 7972 5400
rect 7005 5342 7972 5344
rect 7005 5339 7071 5342
rect 7966 5340 7972 5342
rect 8036 5402 8042 5404
rect 8477 5402 8543 5405
rect 8036 5400 8543 5402
rect 8036 5344 8482 5400
rect 8538 5344 8543 5400
rect 8036 5342 8543 5344
rect 8036 5340 8042 5342
rect 8477 5339 8543 5342
rect 9254 5340 9260 5404
rect 9324 5402 9330 5404
rect 11700 5402 11760 5478
rect 11881 5475 11947 5478
rect 12022 5478 12204 5538
rect 9324 5342 11760 5402
rect 11881 5402 11947 5405
rect 12022 5402 12082 5478
rect 12198 5476 12204 5478
rect 12268 5476 12274 5540
rect 12790 5472 13106 5473
rect 12790 5408 12796 5472
rect 12860 5408 12876 5472
rect 12940 5408 12956 5472
rect 13020 5408 13036 5472
rect 13100 5408 13106 5472
rect 12790 5407 13106 5408
rect 11881 5400 12082 5402
rect 11881 5344 11886 5400
rect 11942 5344 12082 5400
rect 11881 5342 12082 5344
rect 12157 5402 12223 5405
rect 12525 5402 12591 5405
rect 12157 5400 12591 5402
rect 12157 5344 12162 5400
rect 12218 5344 12530 5400
rect 12586 5344 12591 5400
rect 12157 5342 12591 5344
rect 9324 5340 9330 5342
rect 11881 5339 11947 5342
rect 12157 5339 12223 5342
rect 12525 5339 12591 5342
rect 0 5266 400 5296
rect 2773 5266 2839 5269
rect 0 5264 2839 5266
rect 0 5208 2778 5264
rect 2834 5208 2839 5264
rect 0 5206 2839 5208
rect 0 5176 400 5206
rect 2773 5203 2839 5206
rect 6678 5204 6684 5268
rect 6748 5266 6754 5268
rect 9489 5266 9555 5269
rect 9765 5266 9831 5269
rect 15745 5266 15811 5269
rect 6748 5264 15811 5266
rect 6748 5208 9494 5264
rect 9550 5208 9770 5264
rect 9826 5208 15750 5264
rect 15806 5208 15811 5264
rect 6748 5206 15811 5208
rect 6748 5204 6754 5206
rect 9489 5203 9555 5206
rect 9765 5203 9831 5206
rect 15745 5203 15811 5206
rect 5165 5130 5231 5133
rect 6126 5130 6132 5132
rect 5165 5128 6132 5130
rect 5165 5072 5170 5128
rect 5226 5072 6132 5128
rect 5165 5070 6132 5072
rect 5165 5067 5231 5070
rect 6126 5068 6132 5070
rect 6196 5068 6202 5132
rect 6637 5130 6703 5133
rect 8017 5130 8083 5133
rect 8753 5130 8819 5133
rect 9581 5130 9647 5133
rect 12157 5130 12223 5133
rect 6637 5128 7344 5130
rect 6637 5072 6642 5128
rect 6698 5072 7344 5128
rect 6637 5070 7344 5072
rect 6637 5067 6703 5070
rect 3325 4994 3391 4997
rect 6640 4994 6700 5067
rect 3325 4992 6700 4994
rect 3325 4936 3330 4992
rect 3386 4936 6700 4992
rect 3325 4934 6700 4936
rect 7284 4994 7344 5070
rect 8017 5128 9647 5130
rect 8017 5072 8022 5128
rect 8078 5072 8758 5128
rect 8814 5072 9586 5128
rect 9642 5072 9647 5128
rect 8017 5070 9647 5072
rect 8017 5067 8083 5070
rect 8753 5067 8819 5070
rect 9581 5067 9647 5070
rect 10366 5128 12223 5130
rect 10366 5072 12162 5128
rect 12218 5072 12223 5128
rect 10366 5070 12223 5072
rect 10366 4996 10426 5070
rect 12157 5067 12223 5070
rect 12341 5130 12407 5133
rect 14457 5130 14523 5133
rect 12341 5128 14523 5130
rect 12341 5072 12346 5128
rect 12402 5072 14462 5128
rect 14518 5072 14523 5128
rect 12341 5070 14523 5072
rect 12341 5067 12407 5070
rect 14457 5067 14523 5070
rect 15142 5068 15148 5132
rect 15212 5130 15218 5132
rect 15285 5130 15351 5133
rect 15212 5128 15351 5130
rect 15212 5072 15290 5128
rect 15346 5072 15351 5128
rect 15212 5070 15351 5072
rect 15212 5068 15218 5070
rect 15285 5067 15351 5070
rect 10358 4994 10364 4996
rect 7284 4934 10364 4994
rect 3325 4931 3391 4934
rect 10358 4932 10364 4934
rect 10428 4932 10434 4996
rect 11605 4994 11671 4997
rect 12014 4994 12020 4996
rect 11605 4992 12020 4994
rect 11605 4936 11610 4992
rect 11666 4936 12020 4992
rect 11605 4934 12020 4936
rect 11605 4931 11671 4934
rect 12014 4932 12020 4934
rect 12084 4932 12090 4996
rect 12198 4932 12204 4996
rect 12268 4994 12274 4996
rect 12617 4994 12683 4997
rect 12268 4992 12683 4994
rect 12268 4936 12622 4992
rect 12678 4936 12683 4992
rect 12268 4934 12683 4936
rect 12268 4932 12274 4934
rect 12617 4931 12683 4934
rect 2920 4928 3236 4929
rect 2920 4864 2926 4928
rect 2990 4864 3006 4928
rect 3070 4864 3086 4928
rect 3150 4864 3166 4928
rect 3230 4864 3236 4928
rect 2920 4863 3236 4864
rect 6868 4928 7184 4929
rect 6868 4864 6874 4928
rect 6938 4864 6954 4928
rect 7018 4864 7034 4928
rect 7098 4864 7114 4928
rect 7178 4864 7184 4928
rect 6868 4863 7184 4864
rect 10816 4928 11132 4929
rect 10816 4864 10822 4928
rect 10886 4864 10902 4928
rect 10966 4864 10982 4928
rect 11046 4864 11062 4928
rect 11126 4864 11132 4928
rect 10816 4863 11132 4864
rect 14764 4928 15080 4929
rect 14764 4864 14770 4928
rect 14834 4864 14850 4928
rect 14914 4864 14930 4928
rect 14994 4864 15010 4928
rect 15074 4864 15080 4928
rect 14764 4863 15080 4864
rect 8702 4796 8708 4860
rect 8772 4858 8778 4860
rect 8845 4858 8911 4861
rect 9673 4858 9739 4861
rect 8772 4856 9739 4858
rect 8772 4800 8850 4856
rect 8906 4800 9678 4856
rect 9734 4800 9739 4856
rect 8772 4798 9739 4800
rect 8772 4796 8778 4798
rect 8845 4795 8911 4798
rect 9673 4795 9739 4798
rect 9806 4796 9812 4860
rect 9876 4858 9882 4860
rect 10593 4858 10659 4861
rect 9876 4856 10659 4858
rect 9876 4800 10598 4856
rect 10654 4800 10659 4856
rect 9876 4798 10659 4800
rect 9876 4796 9882 4798
rect 10593 4795 10659 4798
rect 11830 4796 11836 4860
rect 11900 4858 11906 4860
rect 12801 4858 12867 4861
rect 11900 4856 12867 4858
rect 11900 4800 12806 4856
rect 12862 4800 12867 4856
rect 11900 4798 12867 4800
rect 11900 4796 11906 4798
rect 2497 4722 2563 4725
rect 6637 4722 6703 4725
rect 2497 4720 6703 4722
rect 2497 4664 2502 4720
rect 2558 4664 6642 4720
rect 6698 4664 6703 4720
rect 2497 4662 6703 4664
rect 2497 4659 2563 4662
rect 6637 4659 6703 4662
rect 6913 4722 6979 4725
rect 9673 4724 9739 4725
rect 9622 4722 9628 4724
rect 6913 4720 9460 4722
rect 6913 4664 6918 4720
rect 6974 4664 9460 4720
rect 6913 4662 9460 4664
rect 9582 4662 9628 4722
rect 9692 4720 9739 4724
rect 9734 4664 9739 4720
rect 6913 4659 6979 4662
rect 3785 4586 3851 4589
rect 5533 4586 5599 4589
rect 3785 4584 5599 4586
rect 3785 4528 3790 4584
rect 3846 4528 5538 4584
rect 5594 4528 5599 4584
rect 3785 4526 5599 4528
rect 3785 4523 3851 4526
rect 5533 4523 5599 4526
rect 6821 4586 6887 4589
rect 7782 4586 7788 4588
rect 6821 4584 7788 4586
rect 6821 4528 6826 4584
rect 6882 4528 7788 4584
rect 6821 4526 7788 4528
rect 6821 4523 6887 4526
rect 7782 4524 7788 4526
rect 7852 4524 7858 4588
rect 8293 4586 8359 4589
rect 9400 4586 9460 4662
rect 9622 4660 9628 4662
rect 9692 4660 9739 4664
rect 9806 4660 9812 4724
rect 9876 4722 9882 4724
rect 10225 4722 10291 4725
rect 11278 4722 11284 4724
rect 9876 4720 11284 4722
rect 9876 4664 10230 4720
rect 10286 4664 11284 4720
rect 9876 4662 11284 4664
rect 9876 4660 9882 4662
rect 9673 4659 9739 4660
rect 10225 4659 10291 4662
rect 11278 4660 11284 4662
rect 11348 4660 11354 4724
rect 11838 4586 11898 4796
rect 12801 4795 12867 4798
rect 13486 4796 13492 4860
rect 13556 4858 13562 4860
rect 14273 4858 14339 4861
rect 13556 4856 14339 4858
rect 13556 4800 14278 4856
rect 14334 4800 14339 4856
rect 13556 4798 14339 4800
rect 13556 4796 13562 4798
rect 14273 4795 14339 4798
rect 12014 4660 12020 4724
rect 12084 4722 12090 4724
rect 13302 4722 13308 4724
rect 12084 4662 13308 4722
rect 12084 4660 12090 4662
rect 13302 4660 13308 4662
rect 13372 4660 13378 4724
rect 8293 4584 9322 4586
rect 8293 4528 8298 4584
rect 8354 4528 9322 4584
rect 8293 4526 9322 4528
rect 9400 4526 11898 4586
rect 11973 4586 12039 4589
rect 13537 4586 13603 4589
rect 11973 4584 13603 4586
rect 11973 4528 11978 4584
rect 12034 4528 13542 4584
rect 13598 4528 13603 4584
rect 11973 4526 13603 4528
rect 8293 4523 8359 4526
rect 5809 4450 5875 4453
rect 7373 4450 7439 4453
rect 9262 4450 9322 4526
rect 11973 4523 12039 4526
rect 13537 4523 13603 4526
rect 12065 4450 12131 4453
rect 5809 4448 7252 4450
rect 5809 4392 5814 4448
rect 5870 4392 7252 4448
rect 5809 4390 7252 4392
rect 5809 4387 5875 4390
rect 4894 4384 5210 4385
rect 4894 4320 4900 4384
rect 4964 4320 4980 4384
rect 5044 4320 5060 4384
rect 5124 4320 5140 4384
rect 5204 4320 5210 4384
rect 4894 4319 5210 4320
rect 2865 4314 2931 4317
rect 3601 4314 3667 4317
rect 2865 4312 3667 4314
rect 2865 4256 2870 4312
rect 2926 4256 3606 4312
rect 3662 4256 3667 4312
rect 2865 4254 3667 4256
rect 7192 4314 7252 4390
rect 7373 4448 8218 4450
rect 7373 4392 7378 4448
rect 7434 4392 8218 4448
rect 7373 4390 8218 4392
rect 9262 4448 12131 4450
rect 9262 4392 12070 4448
rect 12126 4392 12131 4448
rect 9262 4390 12131 4392
rect 7373 4387 7439 4390
rect 8017 4314 8083 4317
rect 7192 4312 8083 4314
rect 7192 4256 8022 4312
rect 8078 4256 8083 4312
rect 7192 4254 8083 4256
rect 8158 4314 8218 4390
rect 12065 4387 12131 4390
rect 14222 4388 14228 4452
rect 14292 4450 14298 4452
rect 14641 4450 14707 4453
rect 14292 4448 14707 4450
rect 14292 4392 14646 4448
rect 14702 4392 14707 4448
rect 14292 4390 14707 4392
rect 14292 4388 14298 4390
rect 14641 4387 14707 4390
rect 8842 4384 9158 4385
rect 8842 4320 8848 4384
rect 8912 4320 8928 4384
rect 8992 4320 9008 4384
rect 9072 4320 9088 4384
rect 9152 4320 9158 4384
rect 8842 4319 9158 4320
rect 12790 4384 13106 4385
rect 12790 4320 12796 4384
rect 12860 4320 12876 4384
rect 12940 4320 12956 4384
rect 13020 4320 13036 4384
rect 13100 4320 13106 4384
rect 12790 4319 13106 4320
rect 8702 4314 8708 4316
rect 8158 4254 8708 4314
rect 2865 4251 2931 4254
rect 3601 4251 3667 4254
rect 8017 4251 8083 4254
rect 8702 4252 8708 4254
rect 8772 4252 8778 4316
rect 9305 4314 9371 4317
rect 10685 4314 10751 4317
rect 9305 4312 10751 4314
rect 9305 4256 9310 4312
rect 9366 4256 10690 4312
rect 10746 4256 10751 4312
rect 9305 4254 10751 4256
rect 9305 4251 9371 4254
rect 10685 4251 10751 4254
rect 11237 4314 11303 4317
rect 11881 4314 11947 4317
rect 12617 4314 12683 4317
rect 11237 4312 11947 4314
rect 11237 4256 11242 4312
rect 11298 4256 11886 4312
rect 11942 4256 11947 4312
rect 11237 4254 11947 4256
rect 11237 4251 11303 4254
rect 11881 4251 11947 4254
rect 12206 4312 12683 4314
rect 12206 4256 12622 4312
rect 12678 4256 12683 4312
rect 12206 4254 12683 4256
rect 7966 4116 7972 4180
rect 8036 4178 8042 4180
rect 12206 4178 12266 4254
rect 12617 4251 12683 4254
rect 14089 4314 14155 4317
rect 17217 4314 17283 4317
rect 14089 4312 17283 4314
rect 14089 4256 14094 4312
rect 14150 4256 17222 4312
rect 17278 4256 17283 4312
rect 14089 4254 17283 4256
rect 14089 4251 14155 4254
rect 17217 4251 17283 4254
rect 8036 4118 12266 4178
rect 12341 4178 12407 4181
rect 15510 4178 15516 4180
rect 12341 4176 15516 4178
rect 12341 4120 12346 4176
rect 12402 4120 15516 4176
rect 12341 4118 15516 4120
rect 8036 4116 8042 4118
rect 12341 4115 12407 4118
rect 15510 4116 15516 4118
rect 15580 4116 15586 4180
rect 16021 4178 16087 4181
rect 16798 4178 16804 4180
rect 16021 4176 16804 4178
rect 16021 4120 16026 4176
rect 16082 4120 16804 4176
rect 16021 4118 16804 4120
rect 16021 4115 16087 4118
rect 16798 4116 16804 4118
rect 16868 4116 16874 4180
rect 4797 4042 4863 4045
rect 13721 4042 13787 4045
rect 15009 4042 15075 4045
rect 4797 4040 13787 4042
rect 4797 3984 4802 4040
rect 4858 3984 13726 4040
rect 13782 3984 13787 4040
rect 4797 3982 13787 3984
rect 4797 3979 4863 3982
rect 13721 3979 13787 3982
rect 14368 4040 15075 4042
rect 14368 3984 15014 4040
rect 15070 3984 15075 4040
rect 14368 3982 15075 3984
rect 14368 3909 14428 3982
rect 15009 3979 15075 3982
rect 4429 3906 4495 3909
rect 6310 3906 6316 3908
rect 4429 3904 6316 3906
rect 4429 3848 4434 3904
rect 4490 3848 6316 3904
rect 4429 3846 6316 3848
rect 4429 3843 4495 3846
rect 6310 3844 6316 3846
rect 6380 3844 6386 3908
rect 6453 3906 6519 3909
rect 6637 3906 6703 3909
rect 7373 3908 7439 3909
rect 7373 3906 7420 3908
rect 6453 3904 6703 3906
rect 6453 3848 6458 3904
rect 6514 3848 6642 3904
rect 6698 3848 6703 3904
rect 6453 3846 6703 3848
rect 7328 3904 7420 3906
rect 7328 3848 7378 3904
rect 7328 3846 7420 3848
rect 6453 3843 6519 3846
rect 6637 3843 6703 3846
rect 7373 3844 7420 3846
rect 7484 3844 7490 3908
rect 7782 3844 7788 3908
rect 7852 3906 7858 3908
rect 9990 3906 9996 3908
rect 7852 3846 9996 3906
rect 7852 3844 7858 3846
rect 9990 3844 9996 3846
rect 10060 3906 10066 3908
rect 10501 3906 10567 3909
rect 10060 3904 10567 3906
rect 10060 3848 10506 3904
rect 10562 3848 10567 3904
rect 10060 3846 10567 3848
rect 10060 3844 10066 3846
rect 7373 3843 7439 3844
rect 10501 3843 10567 3846
rect 11237 3906 11303 3909
rect 12014 3906 12020 3908
rect 11237 3904 12020 3906
rect 11237 3848 11242 3904
rect 11298 3848 12020 3904
rect 11237 3846 12020 3848
rect 11237 3843 11303 3846
rect 12014 3844 12020 3846
rect 12084 3844 12090 3908
rect 12617 3906 12683 3909
rect 13169 3906 13235 3909
rect 12617 3904 13235 3906
rect 12617 3848 12622 3904
rect 12678 3848 13174 3904
rect 13230 3848 13235 3904
rect 12617 3846 13235 3848
rect 12617 3843 12683 3846
rect 13169 3843 13235 3846
rect 13721 3906 13787 3909
rect 14089 3906 14155 3909
rect 13721 3904 14155 3906
rect 13721 3848 13726 3904
rect 13782 3848 14094 3904
rect 14150 3848 14155 3904
rect 13721 3846 14155 3848
rect 13721 3843 13787 3846
rect 14089 3843 14155 3846
rect 14365 3904 14431 3909
rect 14365 3848 14370 3904
rect 14426 3848 14431 3904
rect 14365 3843 14431 3848
rect 2920 3840 3236 3841
rect 0 3770 400 3800
rect 2920 3776 2926 3840
rect 2990 3776 3006 3840
rect 3070 3776 3086 3840
rect 3150 3776 3166 3840
rect 3230 3776 3236 3840
rect 2920 3775 3236 3776
rect 6868 3840 7184 3841
rect 6868 3776 6874 3840
rect 6938 3776 6954 3840
rect 7018 3776 7034 3840
rect 7098 3776 7114 3840
rect 7178 3776 7184 3840
rect 6868 3775 7184 3776
rect 10816 3840 11132 3841
rect 10816 3776 10822 3840
rect 10886 3776 10902 3840
rect 10966 3776 10982 3840
rect 11046 3776 11062 3840
rect 11126 3776 11132 3840
rect 10816 3775 11132 3776
rect 14764 3840 15080 3841
rect 14764 3776 14770 3840
rect 14834 3776 14850 3840
rect 14914 3776 14930 3840
rect 14994 3776 15010 3840
rect 15074 3776 15080 3840
rect 14764 3775 15080 3776
rect 5809 3772 5875 3773
rect 0 3710 2790 3770
rect 0 3680 400 3710
rect 2730 3634 2790 3710
rect 5758 3708 5764 3772
rect 5828 3770 5875 3772
rect 8017 3770 8083 3773
rect 8334 3770 8340 3772
rect 5828 3768 5920 3770
rect 5870 3712 5920 3768
rect 5828 3710 5920 3712
rect 8017 3768 8340 3770
rect 8017 3712 8022 3768
rect 8078 3712 8340 3768
rect 8017 3710 8340 3712
rect 5828 3708 5875 3710
rect 5809 3707 5875 3708
rect 8017 3707 8083 3710
rect 8334 3708 8340 3710
rect 8404 3708 8410 3772
rect 8702 3708 8708 3772
rect 8772 3770 8778 3772
rect 9121 3770 9187 3773
rect 8772 3768 9187 3770
rect 8772 3712 9126 3768
rect 9182 3712 9187 3768
rect 8772 3710 9187 3712
rect 8772 3708 8778 3710
rect 9121 3707 9187 3710
rect 11646 3708 11652 3772
rect 11716 3770 11722 3772
rect 12801 3770 12867 3773
rect 11716 3768 12867 3770
rect 11716 3712 12806 3768
rect 12862 3712 12867 3768
rect 11716 3710 12867 3712
rect 11716 3708 11722 3710
rect 12801 3707 12867 3710
rect 3693 3634 3759 3637
rect 2730 3632 3759 3634
rect 2730 3576 3698 3632
rect 3754 3576 3759 3632
rect 2730 3574 3759 3576
rect 3693 3571 3759 3574
rect 3877 3634 3943 3637
rect 11697 3634 11763 3637
rect 14038 3634 14044 3636
rect 3877 3632 11763 3634
rect 3877 3576 3882 3632
rect 3938 3576 11702 3632
rect 11758 3576 11763 3632
rect 3877 3574 11763 3576
rect 3877 3571 3943 3574
rect 11697 3571 11763 3574
rect 11838 3574 14044 3634
rect 2630 3436 2636 3500
rect 2700 3498 2706 3500
rect 3141 3498 3207 3501
rect 2700 3496 3207 3498
rect 2700 3440 3146 3496
rect 3202 3440 3207 3496
rect 2700 3438 3207 3440
rect 2700 3436 2706 3438
rect 3141 3435 3207 3438
rect 5993 3498 6059 3501
rect 8017 3500 8083 3501
rect 7966 3498 7972 3500
rect 5993 3496 7972 3498
rect 8036 3496 8083 3500
rect 5993 3440 5998 3496
rect 6054 3440 7972 3496
rect 8078 3440 8083 3496
rect 5993 3438 7972 3440
rect 5993 3435 6059 3438
rect 7966 3436 7972 3438
rect 8036 3436 8083 3440
rect 8017 3435 8083 3436
rect 8477 3498 8543 3501
rect 11838 3498 11898 3574
rect 14038 3572 14044 3574
rect 14108 3572 14114 3636
rect 8477 3496 11898 3498
rect 8477 3440 8482 3496
rect 8538 3440 11898 3496
rect 8477 3438 11898 3440
rect 12801 3498 12867 3501
rect 14549 3498 14615 3501
rect 12801 3496 14615 3498
rect 12801 3440 12806 3496
rect 12862 3440 14554 3496
rect 14610 3440 14615 3496
rect 12801 3438 14615 3440
rect 8477 3435 8543 3438
rect 12801 3435 12867 3438
rect 14549 3435 14615 3438
rect 4153 3362 4219 3365
rect 4286 3362 4292 3364
rect 4153 3360 4292 3362
rect 4153 3304 4158 3360
rect 4214 3304 4292 3360
rect 4153 3302 4292 3304
rect 4153 3299 4219 3302
rect 4286 3300 4292 3302
rect 4356 3300 4362 3364
rect 7005 3362 7071 3365
rect 7598 3362 7604 3364
rect 7005 3360 7604 3362
rect 7005 3304 7010 3360
rect 7066 3304 7604 3360
rect 7005 3302 7604 3304
rect 7005 3299 7071 3302
rect 7598 3300 7604 3302
rect 7668 3300 7674 3364
rect 8201 3362 8267 3365
rect 8518 3362 8524 3364
rect 8201 3360 8524 3362
rect 8201 3304 8206 3360
rect 8262 3304 8524 3360
rect 8201 3302 8524 3304
rect 8201 3299 8267 3302
rect 8518 3300 8524 3302
rect 8588 3300 8594 3364
rect 9305 3362 9371 3365
rect 11881 3362 11947 3365
rect 9305 3360 11947 3362
rect 9305 3304 9310 3360
rect 9366 3304 11886 3360
rect 11942 3304 11947 3360
rect 9305 3302 11947 3304
rect 9305 3299 9371 3302
rect 11881 3299 11947 3302
rect 13721 3362 13787 3365
rect 17585 3362 17651 3365
rect 13721 3360 17651 3362
rect 13721 3304 13726 3360
rect 13782 3304 17590 3360
rect 17646 3304 17651 3360
rect 13721 3302 17651 3304
rect 13721 3299 13787 3302
rect 17585 3299 17651 3302
rect 4894 3296 5210 3297
rect 4894 3232 4900 3296
rect 4964 3232 4980 3296
rect 5044 3232 5060 3296
rect 5124 3232 5140 3296
rect 5204 3232 5210 3296
rect 4894 3231 5210 3232
rect 1485 3226 1551 3229
rect 5441 3226 5507 3229
rect 5574 3226 5580 3228
rect 1485 3224 4722 3226
rect 1485 3168 1490 3224
rect 1546 3168 4722 3224
rect 1485 3166 4722 3168
rect 1485 3163 1551 3166
rect 4662 3090 4722 3166
rect 5441 3224 5580 3226
rect 5441 3168 5446 3224
rect 5502 3168 5580 3224
rect 5441 3166 5580 3168
rect 5441 3163 5507 3166
rect 5574 3164 5580 3166
rect 5644 3164 5650 3228
rect 6545 3226 6611 3229
rect 8204 3226 8264 3299
rect 8842 3296 9158 3297
rect 8842 3232 8848 3296
rect 8912 3232 8928 3296
rect 8992 3232 9008 3296
rect 9072 3232 9088 3296
rect 9152 3232 9158 3296
rect 8842 3231 9158 3232
rect 12790 3296 13106 3297
rect 12790 3232 12796 3296
rect 12860 3232 12876 3296
rect 12940 3232 12956 3296
rect 13020 3232 13036 3296
rect 13100 3232 13106 3296
rect 12790 3231 13106 3232
rect 9305 3228 9371 3229
rect 6545 3224 8264 3226
rect 6545 3168 6550 3224
rect 6606 3168 8264 3224
rect 6545 3166 8264 3168
rect 6545 3163 6611 3166
rect 9254 3164 9260 3228
rect 9324 3226 9371 3228
rect 10225 3226 10291 3229
rect 12617 3226 12683 3229
rect 15653 3226 15719 3229
rect 9324 3224 9416 3226
rect 9366 3168 9416 3224
rect 9324 3166 9416 3168
rect 10225 3224 12683 3226
rect 10225 3168 10230 3224
rect 10286 3168 12622 3224
rect 12678 3168 12683 3224
rect 10225 3166 12683 3168
rect 9324 3164 9371 3166
rect 9305 3163 9371 3164
rect 10225 3163 10291 3166
rect 12617 3163 12683 3166
rect 13172 3224 15719 3226
rect 13172 3168 15658 3224
rect 15714 3168 15719 3224
rect 13172 3166 15719 3168
rect 5993 3090 6059 3093
rect 4662 3088 6059 3090
rect 4662 3032 5998 3088
rect 6054 3032 6059 3088
rect 4662 3030 6059 3032
rect 5993 3027 6059 3030
rect 6177 3090 6243 3093
rect 9397 3090 9463 3093
rect 6177 3088 9463 3090
rect 6177 3032 6182 3088
rect 6238 3032 9402 3088
rect 9458 3032 9463 3088
rect 6177 3030 9463 3032
rect 6177 3027 6243 3030
rect 9397 3027 9463 3030
rect 10542 3028 10548 3092
rect 10612 3090 10618 3092
rect 10961 3090 11027 3093
rect 10612 3088 11027 3090
rect 10612 3032 10966 3088
rect 11022 3032 11027 3088
rect 10612 3030 11027 3032
rect 10612 3028 10618 3030
rect 10961 3027 11027 3030
rect 11697 3090 11763 3093
rect 13172 3090 13232 3166
rect 15653 3163 15719 3166
rect 11697 3088 13232 3090
rect 11697 3032 11702 3088
rect 11758 3032 13232 3088
rect 11697 3030 13232 3032
rect 11697 3027 11763 3030
rect 13486 3028 13492 3092
rect 13556 3090 13562 3092
rect 13721 3090 13787 3093
rect 13556 3088 13787 3090
rect 13556 3032 13726 3088
rect 13782 3032 13787 3088
rect 13556 3030 13787 3032
rect 13556 3028 13562 3030
rect 13721 3027 13787 3030
rect 14089 3090 14155 3093
rect 15745 3090 15811 3093
rect 16062 3090 16068 3092
rect 14089 3088 16068 3090
rect 14089 3032 14094 3088
rect 14150 3032 15750 3088
rect 15806 3032 16068 3088
rect 14089 3030 16068 3032
rect 14089 3027 14155 3030
rect 15745 3027 15811 3030
rect 16062 3028 16068 3030
rect 16132 3028 16138 3092
rect 1025 2954 1091 2957
rect 15285 2954 15351 2957
rect 1025 2952 15351 2954
rect 1025 2896 1030 2952
rect 1086 2896 15290 2952
rect 15346 2896 15351 2952
rect 1025 2894 15351 2896
rect 1025 2891 1091 2894
rect 15285 2891 15351 2894
rect 4102 2756 4108 2820
rect 4172 2818 4178 2820
rect 4429 2818 4495 2821
rect 4172 2816 4495 2818
rect 4172 2760 4434 2816
rect 4490 2760 4495 2816
rect 4172 2758 4495 2760
rect 4172 2756 4178 2758
rect 4429 2755 4495 2758
rect 7281 2818 7347 2821
rect 10225 2818 10291 2821
rect 7281 2816 10291 2818
rect 7281 2760 7286 2816
rect 7342 2760 10230 2816
rect 10286 2760 10291 2816
rect 7281 2758 10291 2760
rect 7281 2755 7347 2758
rect 10225 2755 10291 2758
rect 12382 2756 12388 2820
rect 12452 2818 12458 2820
rect 13537 2818 13603 2821
rect 12452 2816 13603 2818
rect 12452 2760 13542 2816
rect 13598 2760 13603 2816
rect 12452 2758 13603 2760
rect 12452 2756 12458 2758
rect 13537 2755 13603 2758
rect 2920 2752 3236 2753
rect 2920 2688 2926 2752
rect 2990 2688 3006 2752
rect 3070 2688 3086 2752
rect 3150 2688 3166 2752
rect 3230 2688 3236 2752
rect 2920 2687 3236 2688
rect 6868 2752 7184 2753
rect 6868 2688 6874 2752
rect 6938 2688 6954 2752
rect 7018 2688 7034 2752
rect 7098 2688 7114 2752
rect 7178 2688 7184 2752
rect 6868 2687 7184 2688
rect 10816 2752 11132 2753
rect 10816 2688 10822 2752
rect 10886 2688 10902 2752
rect 10966 2688 10982 2752
rect 11046 2688 11062 2752
rect 11126 2688 11132 2752
rect 10816 2687 11132 2688
rect 14764 2752 15080 2753
rect 14764 2688 14770 2752
rect 14834 2688 14850 2752
rect 14914 2688 14930 2752
rect 14994 2688 15010 2752
rect 15074 2688 15080 2752
rect 14764 2687 15080 2688
rect 7557 2682 7623 2685
rect 10174 2682 10180 2684
rect 7557 2680 10180 2682
rect 7557 2624 7562 2680
rect 7618 2624 10180 2680
rect 7557 2622 10180 2624
rect 7557 2619 7623 2622
rect 10174 2620 10180 2622
rect 10244 2620 10250 2684
rect 12065 2682 12131 2685
rect 12198 2682 12204 2684
rect 12065 2680 12204 2682
rect 12065 2624 12070 2680
rect 12126 2624 12204 2680
rect 12065 2622 12204 2624
rect 12065 2619 12131 2622
rect 12198 2620 12204 2622
rect 12268 2620 12274 2684
rect 12341 2682 12407 2685
rect 13997 2682 14063 2685
rect 12341 2680 14063 2682
rect 12341 2624 12346 2680
rect 12402 2624 14002 2680
rect 14058 2624 14063 2680
rect 12341 2622 14063 2624
rect 12341 2619 12407 2622
rect 13997 2619 14063 2622
rect 13 2546 79 2549
rect 2865 2546 2931 2549
rect 6637 2546 6703 2549
rect 8201 2546 8267 2549
rect 9806 2546 9812 2548
rect 13 2544 536 2546
rect 13 2488 18 2544
rect 74 2488 536 2544
rect 13 2486 536 2488
rect 13 2483 79 2486
rect 0 2274 400 2304
rect 476 2274 536 2486
rect 2865 2544 6703 2546
rect 2865 2488 2870 2544
rect 2926 2488 6642 2544
rect 6698 2488 6703 2544
rect 2865 2486 6703 2488
rect 2865 2483 2931 2486
rect 6637 2483 6703 2486
rect 6824 2544 8267 2546
rect 6824 2488 8206 2544
rect 8262 2488 8267 2544
rect 6824 2486 8267 2488
rect 2497 2410 2563 2413
rect 3141 2410 3207 2413
rect 2497 2408 3207 2410
rect 2497 2352 2502 2408
rect 2558 2352 3146 2408
rect 3202 2352 3207 2408
rect 2497 2350 3207 2352
rect 2497 2347 2563 2350
rect 3141 2347 3207 2350
rect 4153 2410 4219 2413
rect 6824 2410 6884 2486
rect 8201 2483 8267 2486
rect 8572 2486 9812 2546
rect 4153 2408 6884 2410
rect 4153 2352 4158 2408
rect 4214 2352 6884 2408
rect 4153 2350 6884 2352
rect 7649 2410 7715 2413
rect 8572 2410 8632 2486
rect 9806 2484 9812 2486
rect 9876 2484 9882 2548
rect 10869 2546 10935 2549
rect 16021 2546 16087 2549
rect 10869 2544 16087 2546
rect 10869 2488 10874 2544
rect 10930 2488 16026 2544
rect 16082 2488 16087 2544
rect 10869 2486 16087 2488
rect 10869 2483 10935 2486
rect 16021 2483 16087 2486
rect 7649 2408 8632 2410
rect 7649 2352 7654 2408
rect 7710 2352 8632 2408
rect 7649 2350 8632 2352
rect 8753 2410 8819 2413
rect 12157 2410 12223 2413
rect 14641 2410 14707 2413
rect 8753 2408 12223 2410
rect 8753 2352 8758 2408
rect 8814 2352 12162 2408
rect 12218 2352 12223 2408
rect 8753 2350 12223 2352
rect 4153 2347 4219 2350
rect 7649 2347 7715 2350
rect 8753 2347 8819 2350
rect 12157 2347 12223 2350
rect 12390 2408 14707 2410
rect 12390 2352 14646 2408
rect 14702 2352 14707 2408
rect 12390 2350 14707 2352
rect 0 2214 536 2274
rect 5993 2274 6059 2277
rect 7782 2274 7788 2276
rect 5993 2272 7788 2274
rect 5993 2216 5998 2272
rect 6054 2216 7788 2272
rect 5993 2214 7788 2216
rect 0 2184 400 2214
rect 5993 2211 6059 2214
rect 7782 2212 7788 2214
rect 7852 2212 7858 2276
rect 8150 2212 8156 2276
rect 8220 2274 8226 2276
rect 8385 2274 8451 2277
rect 8220 2272 8451 2274
rect 8220 2216 8390 2272
rect 8446 2216 8451 2272
rect 8220 2214 8451 2216
rect 8220 2212 8226 2214
rect 8385 2211 8451 2214
rect 9305 2274 9371 2277
rect 12390 2274 12450 2350
rect 14641 2347 14707 2350
rect 15009 2410 15075 2413
rect 15326 2410 15332 2412
rect 15009 2408 15332 2410
rect 15009 2352 15014 2408
rect 15070 2352 15332 2408
rect 15009 2350 15332 2352
rect 15009 2347 15075 2350
rect 15326 2348 15332 2350
rect 15396 2348 15402 2412
rect 9305 2272 12450 2274
rect 9305 2216 9310 2272
rect 9366 2216 12450 2272
rect 9305 2214 12450 2216
rect 13169 2272 13235 2277
rect 13169 2216 13174 2272
rect 13230 2216 13235 2272
rect 9305 2211 9371 2214
rect 13169 2211 13235 2216
rect 4894 2208 5210 2209
rect 4894 2144 4900 2208
rect 4964 2144 4980 2208
rect 5044 2144 5060 2208
rect 5124 2144 5140 2208
rect 5204 2144 5210 2208
rect 4894 2143 5210 2144
rect 8842 2208 9158 2209
rect 8842 2144 8848 2208
rect 8912 2144 8928 2208
rect 8992 2144 9008 2208
rect 9072 2144 9088 2208
rect 9152 2144 9158 2208
rect 8842 2143 9158 2144
rect 12790 2208 13106 2209
rect 12790 2144 12796 2208
rect 12860 2144 12876 2208
rect 12940 2144 12956 2208
rect 13020 2144 13036 2208
rect 13100 2144 13106 2208
rect 12790 2143 13106 2144
rect 6085 2138 6151 2141
rect 8201 2138 8267 2141
rect 6085 2136 8267 2138
rect 6085 2080 6090 2136
rect 6146 2080 8206 2136
rect 8262 2080 8267 2136
rect 6085 2078 8267 2080
rect 6085 2075 6151 2078
rect 8201 2075 8267 2078
rect 9438 2076 9444 2140
rect 9508 2138 9514 2140
rect 9857 2138 9923 2141
rect 9508 2136 9923 2138
rect 9508 2080 9862 2136
rect 9918 2080 9923 2136
rect 9508 2078 9923 2080
rect 9508 2076 9514 2078
rect 9857 2075 9923 2078
rect 10358 2076 10364 2140
rect 10428 2138 10434 2140
rect 10777 2138 10843 2141
rect 12433 2140 12499 2141
rect 10428 2136 10843 2138
rect 10428 2080 10782 2136
rect 10838 2080 10843 2136
rect 10428 2078 10843 2080
rect 10428 2076 10434 2078
rect 10777 2075 10843 2078
rect 12382 2076 12388 2140
rect 12452 2138 12499 2140
rect 13172 2138 13232 2211
rect 14825 2138 14891 2141
rect 12452 2136 12544 2138
rect 12494 2080 12544 2136
rect 12452 2078 12544 2080
rect 13172 2136 14891 2138
rect 13172 2080 14830 2136
rect 14886 2080 14891 2136
rect 13172 2078 14891 2080
rect 12452 2076 12499 2078
rect 12433 2075 12499 2076
rect 14825 2075 14891 2078
rect 14549 2002 14615 2005
rect 2730 2000 14615 2002
rect 2730 1944 14554 2000
rect 14610 1944 14615 2000
rect 2730 1942 14615 1944
rect 2730 1869 2790 1942
rect 14549 1939 14615 1942
rect 2681 1864 2790 1869
rect 2681 1808 2686 1864
rect 2742 1808 2790 1864
rect 2681 1806 2790 1808
rect 5165 1866 5231 1869
rect 10133 1866 10199 1869
rect 10869 1866 10935 1869
rect 11789 1866 11855 1869
rect 5165 1864 10199 1866
rect 5165 1808 5170 1864
rect 5226 1808 10138 1864
rect 10194 1808 10199 1864
rect 5165 1806 10199 1808
rect 2681 1803 2747 1806
rect 5165 1803 5231 1806
rect 10133 1803 10199 1806
rect 10688 1864 11855 1866
rect 10688 1808 10874 1864
rect 10930 1808 11794 1864
rect 11850 1808 11855 1864
rect 10688 1806 11855 1808
rect 7833 1730 7899 1733
rect 10688 1730 10748 1806
rect 10869 1803 10935 1806
rect 11789 1803 11855 1806
rect 12985 1866 13051 1869
rect 13670 1866 13676 1868
rect 12985 1864 13676 1866
rect 12985 1808 12990 1864
rect 13046 1808 13676 1864
rect 12985 1806 13676 1808
rect 12985 1803 13051 1806
rect 13670 1804 13676 1806
rect 13740 1804 13746 1868
rect 7833 1728 10748 1730
rect 7833 1672 7838 1728
rect 7894 1672 10748 1728
rect 7833 1670 10748 1672
rect 11329 1730 11395 1733
rect 11462 1730 11468 1732
rect 11329 1728 11468 1730
rect 11329 1672 11334 1728
rect 11390 1672 11468 1728
rect 11329 1670 11468 1672
rect 7833 1667 7899 1670
rect 11329 1667 11395 1670
rect 11462 1668 11468 1670
rect 11532 1668 11538 1732
rect 12566 1668 12572 1732
rect 12636 1730 12642 1732
rect 13261 1730 13327 1733
rect 12636 1728 13327 1730
rect 12636 1672 13266 1728
rect 13322 1672 13327 1728
rect 12636 1670 13327 1672
rect 12636 1668 12642 1670
rect 13261 1667 13327 1670
rect 2920 1664 3236 1665
rect 2920 1600 2926 1664
rect 2990 1600 3006 1664
rect 3070 1600 3086 1664
rect 3150 1600 3166 1664
rect 3230 1600 3236 1664
rect 2920 1599 3236 1600
rect 6868 1664 7184 1665
rect 6868 1600 6874 1664
rect 6938 1600 6954 1664
rect 7018 1600 7034 1664
rect 7098 1600 7114 1664
rect 7178 1600 7184 1664
rect 6868 1599 7184 1600
rect 10816 1664 11132 1665
rect 10816 1600 10822 1664
rect 10886 1600 10902 1664
rect 10966 1600 10982 1664
rect 11046 1600 11062 1664
rect 11126 1600 11132 1664
rect 10816 1599 11132 1600
rect 14764 1664 15080 1665
rect 14764 1600 14770 1664
rect 14834 1600 14850 1664
rect 14914 1600 14930 1664
rect 14994 1600 15010 1664
rect 15074 1600 15080 1664
rect 14764 1599 15080 1600
rect 4061 1594 4127 1597
rect 6269 1594 6335 1597
rect 4061 1592 6335 1594
rect 4061 1536 4066 1592
rect 4122 1536 6274 1592
rect 6330 1536 6335 1592
rect 4061 1534 6335 1536
rect 4061 1531 4127 1534
rect 6269 1531 6335 1534
rect 7281 1594 7347 1597
rect 10225 1594 10291 1597
rect 7281 1592 10291 1594
rect 7281 1536 7286 1592
rect 7342 1536 10230 1592
rect 10286 1536 10291 1592
rect 7281 1534 10291 1536
rect 7281 1531 7347 1534
rect 10225 1531 10291 1534
rect 11697 1594 11763 1597
rect 13486 1594 13492 1596
rect 11697 1592 13492 1594
rect 11697 1536 11702 1592
rect 11758 1536 13492 1592
rect 11697 1534 13492 1536
rect 11697 1531 11763 1534
rect 13486 1532 13492 1534
rect 13556 1532 13562 1596
rect 1301 1458 1367 1461
rect 6821 1458 6887 1461
rect 1301 1456 6887 1458
rect 1301 1400 1306 1456
rect 1362 1400 6826 1456
rect 6882 1400 6887 1456
rect 1301 1398 6887 1400
rect 1301 1395 1367 1398
rect 6821 1395 6887 1398
rect 7005 1458 7071 1461
rect 8150 1458 8156 1460
rect 7005 1456 8156 1458
rect 7005 1400 7010 1456
rect 7066 1400 8156 1456
rect 7005 1398 8156 1400
rect 7005 1395 7071 1398
rect 8150 1396 8156 1398
rect 8220 1396 8226 1460
rect 9213 1458 9279 1461
rect 14365 1458 14431 1461
rect 9213 1456 14431 1458
rect 9213 1400 9218 1456
rect 9274 1400 14370 1456
rect 14426 1400 14431 1456
rect 9213 1398 14431 1400
rect 9213 1395 9279 1398
rect 14365 1395 14431 1398
rect 1485 1322 1551 1325
rect 2957 1322 3023 1325
rect 8753 1322 8819 1325
rect 1485 1320 8819 1322
rect 1485 1264 1490 1320
rect 1546 1264 2962 1320
rect 3018 1264 8758 1320
rect 8814 1264 8819 1320
rect 1485 1262 8819 1264
rect 1485 1259 1551 1262
rect 2957 1259 3023 1262
rect 8753 1259 8819 1262
rect 9949 1322 10015 1325
rect 13537 1322 13603 1325
rect 9949 1320 13603 1322
rect 9949 1264 9954 1320
rect 10010 1264 13542 1320
rect 13598 1264 13603 1320
rect 9949 1262 13603 1264
rect 9949 1259 10015 1262
rect 13537 1259 13603 1262
rect 6453 1186 6519 1189
rect 8569 1186 8635 1189
rect 6453 1184 8635 1186
rect 6453 1128 6458 1184
rect 6514 1128 8574 1184
rect 8630 1128 8635 1184
rect 6453 1126 8635 1128
rect 6453 1123 6519 1126
rect 8569 1123 8635 1126
rect 4894 1120 5210 1121
rect 4894 1056 4900 1120
rect 4964 1056 4980 1120
rect 5044 1056 5060 1120
rect 5124 1056 5140 1120
rect 5204 1056 5210 1120
rect 4894 1055 5210 1056
rect 8842 1120 9158 1121
rect 8842 1056 8848 1120
rect 8912 1056 8928 1120
rect 8992 1056 9008 1120
rect 9072 1056 9088 1120
rect 9152 1056 9158 1120
rect 8842 1055 9158 1056
rect 12790 1120 13106 1121
rect 12790 1056 12796 1120
rect 12860 1056 12876 1120
rect 12940 1056 12956 1120
rect 13020 1056 13036 1120
rect 13100 1056 13106 1120
rect 12790 1055 13106 1056
rect 9489 1050 9555 1053
rect 12525 1050 12591 1053
rect 9489 1048 12591 1050
rect 9489 992 9494 1048
rect 9550 992 12530 1048
rect 12586 992 12591 1048
rect 9489 990 12591 992
rect 9489 987 9555 990
rect 12525 987 12591 990
rect 6177 914 6243 917
rect 14181 914 14247 917
rect 6177 912 14247 914
rect 6177 856 6182 912
rect 6238 856 14186 912
rect 14242 856 14247 912
rect 6177 854 14247 856
rect 6177 851 6243 854
rect 14181 851 14247 854
rect 0 778 400 808
rect 7925 778 7991 781
rect 0 776 7991 778
rect 0 720 7930 776
rect 7986 720 7991 776
rect 0 718 7991 720
rect 0 688 400 718
rect 7925 715 7991 718
rect 8201 778 8267 781
rect 14089 778 14155 781
rect 8201 776 14155 778
rect 8201 720 8206 776
rect 8262 720 14094 776
rect 14150 720 14155 776
rect 8201 718 14155 720
rect 8201 715 8267 718
rect 14089 715 14155 718
rect 1945 642 2011 645
rect 9438 642 9444 644
rect 1945 640 9444 642
rect 1945 584 1950 640
rect 2006 584 9444 640
rect 1945 582 9444 584
rect 1945 579 2011 582
rect 9438 580 9444 582
rect 9508 580 9514 644
rect 11881 642 11947 645
rect 13854 642 13860 644
rect 11881 640 13860 642
rect 11881 584 11886 640
rect 11942 584 13860 640
rect 11881 582 13860 584
rect 11881 579 11947 582
rect 13854 580 13860 582
rect 13924 580 13930 644
rect 9673 506 9739 509
rect 13261 506 13327 509
rect 9673 504 13327 506
rect 9673 448 9678 504
rect 9734 448 13266 504
rect 13322 448 13327 504
rect 9673 446 13327 448
rect 9673 443 9739 446
rect 13261 443 13327 446
<< via3 >>
rect 4900 22876 4964 22880
rect 4900 22820 4904 22876
rect 4904 22820 4960 22876
rect 4960 22820 4964 22876
rect 4900 22816 4964 22820
rect 4980 22876 5044 22880
rect 4980 22820 4984 22876
rect 4984 22820 5040 22876
rect 5040 22820 5044 22876
rect 4980 22816 5044 22820
rect 5060 22876 5124 22880
rect 5060 22820 5064 22876
rect 5064 22820 5120 22876
rect 5120 22820 5124 22876
rect 5060 22816 5124 22820
rect 5140 22876 5204 22880
rect 5140 22820 5144 22876
rect 5144 22820 5200 22876
rect 5200 22820 5204 22876
rect 5140 22816 5204 22820
rect 8848 22876 8912 22880
rect 8848 22820 8852 22876
rect 8852 22820 8908 22876
rect 8908 22820 8912 22876
rect 8848 22816 8912 22820
rect 8928 22876 8992 22880
rect 8928 22820 8932 22876
rect 8932 22820 8988 22876
rect 8988 22820 8992 22876
rect 8928 22816 8992 22820
rect 9008 22876 9072 22880
rect 9008 22820 9012 22876
rect 9012 22820 9068 22876
rect 9068 22820 9072 22876
rect 9008 22816 9072 22820
rect 9088 22876 9152 22880
rect 9088 22820 9092 22876
rect 9092 22820 9148 22876
rect 9148 22820 9152 22876
rect 9088 22816 9152 22820
rect 12796 22876 12860 22880
rect 12796 22820 12800 22876
rect 12800 22820 12856 22876
rect 12856 22820 12860 22876
rect 12796 22816 12860 22820
rect 12876 22876 12940 22880
rect 12876 22820 12880 22876
rect 12880 22820 12936 22876
rect 12936 22820 12940 22876
rect 12876 22816 12940 22820
rect 12956 22876 13020 22880
rect 12956 22820 12960 22876
rect 12960 22820 13016 22876
rect 13016 22820 13020 22876
rect 12956 22816 13020 22820
rect 13036 22876 13100 22880
rect 13036 22820 13040 22876
rect 13040 22820 13096 22876
rect 13096 22820 13100 22876
rect 13036 22816 13100 22820
rect 16620 22476 16684 22540
rect 2926 22332 2990 22336
rect 2926 22276 2930 22332
rect 2930 22276 2986 22332
rect 2986 22276 2990 22332
rect 2926 22272 2990 22276
rect 3006 22332 3070 22336
rect 3006 22276 3010 22332
rect 3010 22276 3066 22332
rect 3066 22276 3070 22332
rect 3006 22272 3070 22276
rect 3086 22332 3150 22336
rect 3086 22276 3090 22332
rect 3090 22276 3146 22332
rect 3146 22276 3150 22332
rect 3086 22272 3150 22276
rect 3166 22332 3230 22336
rect 3166 22276 3170 22332
rect 3170 22276 3226 22332
rect 3226 22276 3230 22332
rect 3166 22272 3230 22276
rect 6874 22332 6938 22336
rect 6874 22276 6878 22332
rect 6878 22276 6934 22332
rect 6934 22276 6938 22332
rect 6874 22272 6938 22276
rect 6954 22332 7018 22336
rect 6954 22276 6958 22332
rect 6958 22276 7014 22332
rect 7014 22276 7018 22332
rect 6954 22272 7018 22276
rect 7034 22332 7098 22336
rect 7034 22276 7038 22332
rect 7038 22276 7094 22332
rect 7094 22276 7098 22332
rect 7034 22272 7098 22276
rect 7114 22332 7178 22336
rect 7114 22276 7118 22332
rect 7118 22276 7174 22332
rect 7174 22276 7178 22332
rect 7114 22272 7178 22276
rect 10822 22332 10886 22336
rect 10822 22276 10826 22332
rect 10826 22276 10882 22332
rect 10882 22276 10886 22332
rect 10822 22272 10886 22276
rect 10902 22332 10966 22336
rect 10902 22276 10906 22332
rect 10906 22276 10962 22332
rect 10962 22276 10966 22332
rect 10902 22272 10966 22276
rect 10982 22332 11046 22336
rect 10982 22276 10986 22332
rect 10986 22276 11042 22332
rect 11042 22276 11046 22332
rect 10982 22272 11046 22276
rect 11062 22332 11126 22336
rect 11062 22276 11066 22332
rect 11066 22276 11122 22332
rect 11122 22276 11126 22332
rect 11062 22272 11126 22276
rect 14770 22332 14834 22336
rect 14770 22276 14774 22332
rect 14774 22276 14830 22332
rect 14830 22276 14834 22332
rect 14770 22272 14834 22276
rect 14850 22332 14914 22336
rect 14850 22276 14854 22332
rect 14854 22276 14910 22332
rect 14910 22276 14914 22332
rect 14850 22272 14914 22276
rect 14930 22332 14994 22336
rect 14930 22276 14934 22332
rect 14934 22276 14990 22332
rect 14990 22276 14994 22332
rect 14930 22272 14994 22276
rect 15010 22332 15074 22336
rect 15010 22276 15014 22332
rect 15014 22276 15070 22332
rect 15070 22276 15074 22332
rect 15010 22272 15074 22276
rect 4900 21788 4964 21792
rect 4900 21732 4904 21788
rect 4904 21732 4960 21788
rect 4960 21732 4964 21788
rect 4900 21728 4964 21732
rect 4980 21788 5044 21792
rect 4980 21732 4984 21788
rect 4984 21732 5040 21788
rect 5040 21732 5044 21788
rect 4980 21728 5044 21732
rect 5060 21788 5124 21792
rect 5060 21732 5064 21788
rect 5064 21732 5120 21788
rect 5120 21732 5124 21788
rect 5060 21728 5124 21732
rect 5140 21788 5204 21792
rect 5140 21732 5144 21788
rect 5144 21732 5200 21788
rect 5200 21732 5204 21788
rect 5140 21728 5204 21732
rect 8848 21788 8912 21792
rect 8848 21732 8852 21788
rect 8852 21732 8908 21788
rect 8908 21732 8912 21788
rect 8848 21728 8912 21732
rect 8928 21788 8992 21792
rect 8928 21732 8932 21788
rect 8932 21732 8988 21788
rect 8988 21732 8992 21788
rect 8928 21728 8992 21732
rect 9008 21788 9072 21792
rect 9008 21732 9012 21788
rect 9012 21732 9068 21788
rect 9068 21732 9072 21788
rect 9008 21728 9072 21732
rect 9088 21788 9152 21792
rect 9088 21732 9092 21788
rect 9092 21732 9148 21788
rect 9148 21732 9152 21788
rect 9088 21728 9152 21732
rect 12796 21788 12860 21792
rect 12796 21732 12800 21788
rect 12800 21732 12856 21788
rect 12856 21732 12860 21788
rect 12796 21728 12860 21732
rect 12876 21788 12940 21792
rect 12876 21732 12880 21788
rect 12880 21732 12936 21788
rect 12936 21732 12940 21788
rect 12876 21728 12940 21732
rect 12956 21788 13020 21792
rect 12956 21732 12960 21788
rect 12960 21732 13016 21788
rect 13016 21732 13020 21788
rect 12956 21728 13020 21732
rect 13036 21788 13100 21792
rect 13036 21732 13040 21788
rect 13040 21732 13096 21788
rect 13096 21732 13100 21788
rect 13036 21728 13100 21732
rect 2926 21244 2990 21248
rect 2926 21188 2930 21244
rect 2930 21188 2986 21244
rect 2986 21188 2990 21244
rect 2926 21184 2990 21188
rect 3006 21244 3070 21248
rect 3006 21188 3010 21244
rect 3010 21188 3066 21244
rect 3066 21188 3070 21244
rect 3006 21184 3070 21188
rect 3086 21244 3150 21248
rect 3086 21188 3090 21244
rect 3090 21188 3146 21244
rect 3146 21188 3150 21244
rect 3086 21184 3150 21188
rect 3166 21244 3230 21248
rect 3166 21188 3170 21244
rect 3170 21188 3226 21244
rect 3226 21188 3230 21244
rect 3166 21184 3230 21188
rect 6874 21244 6938 21248
rect 6874 21188 6878 21244
rect 6878 21188 6934 21244
rect 6934 21188 6938 21244
rect 6874 21184 6938 21188
rect 6954 21244 7018 21248
rect 6954 21188 6958 21244
rect 6958 21188 7014 21244
rect 7014 21188 7018 21244
rect 6954 21184 7018 21188
rect 7034 21244 7098 21248
rect 7034 21188 7038 21244
rect 7038 21188 7094 21244
rect 7094 21188 7098 21244
rect 7034 21184 7098 21188
rect 7114 21244 7178 21248
rect 7114 21188 7118 21244
rect 7118 21188 7174 21244
rect 7174 21188 7178 21244
rect 7114 21184 7178 21188
rect 10822 21244 10886 21248
rect 10822 21188 10826 21244
rect 10826 21188 10882 21244
rect 10882 21188 10886 21244
rect 10822 21184 10886 21188
rect 10902 21244 10966 21248
rect 10902 21188 10906 21244
rect 10906 21188 10962 21244
rect 10962 21188 10966 21244
rect 10902 21184 10966 21188
rect 10982 21244 11046 21248
rect 10982 21188 10986 21244
rect 10986 21188 11042 21244
rect 11042 21188 11046 21244
rect 10982 21184 11046 21188
rect 11062 21244 11126 21248
rect 11062 21188 11066 21244
rect 11066 21188 11122 21244
rect 11122 21188 11126 21244
rect 11062 21184 11126 21188
rect 14770 21244 14834 21248
rect 14770 21188 14774 21244
rect 14774 21188 14830 21244
rect 14830 21188 14834 21244
rect 14770 21184 14834 21188
rect 14850 21244 14914 21248
rect 14850 21188 14854 21244
rect 14854 21188 14910 21244
rect 14910 21188 14914 21244
rect 14850 21184 14914 21188
rect 14930 21244 14994 21248
rect 14930 21188 14934 21244
rect 14934 21188 14990 21244
rect 14990 21188 14994 21244
rect 14930 21184 14994 21188
rect 15010 21244 15074 21248
rect 15010 21188 15014 21244
rect 15014 21188 15070 21244
rect 15070 21188 15074 21244
rect 15010 21184 15074 21188
rect 4900 20700 4964 20704
rect 4900 20644 4904 20700
rect 4904 20644 4960 20700
rect 4960 20644 4964 20700
rect 4900 20640 4964 20644
rect 4980 20700 5044 20704
rect 4980 20644 4984 20700
rect 4984 20644 5040 20700
rect 5040 20644 5044 20700
rect 4980 20640 5044 20644
rect 5060 20700 5124 20704
rect 5060 20644 5064 20700
rect 5064 20644 5120 20700
rect 5120 20644 5124 20700
rect 5060 20640 5124 20644
rect 5140 20700 5204 20704
rect 5140 20644 5144 20700
rect 5144 20644 5200 20700
rect 5200 20644 5204 20700
rect 5140 20640 5204 20644
rect 8848 20700 8912 20704
rect 8848 20644 8852 20700
rect 8852 20644 8908 20700
rect 8908 20644 8912 20700
rect 8848 20640 8912 20644
rect 8928 20700 8992 20704
rect 8928 20644 8932 20700
rect 8932 20644 8988 20700
rect 8988 20644 8992 20700
rect 8928 20640 8992 20644
rect 9008 20700 9072 20704
rect 9008 20644 9012 20700
rect 9012 20644 9068 20700
rect 9068 20644 9072 20700
rect 9008 20640 9072 20644
rect 9088 20700 9152 20704
rect 9088 20644 9092 20700
rect 9092 20644 9148 20700
rect 9148 20644 9152 20700
rect 9088 20640 9152 20644
rect 12796 20700 12860 20704
rect 12796 20644 12800 20700
rect 12800 20644 12856 20700
rect 12856 20644 12860 20700
rect 12796 20640 12860 20644
rect 12876 20700 12940 20704
rect 12876 20644 12880 20700
rect 12880 20644 12936 20700
rect 12936 20644 12940 20700
rect 12876 20640 12940 20644
rect 12956 20700 13020 20704
rect 12956 20644 12960 20700
rect 12960 20644 13016 20700
rect 13016 20644 13020 20700
rect 12956 20640 13020 20644
rect 13036 20700 13100 20704
rect 13036 20644 13040 20700
rect 13040 20644 13096 20700
rect 13096 20644 13100 20700
rect 13036 20640 13100 20644
rect 3740 20300 3804 20364
rect 2926 20156 2990 20160
rect 2926 20100 2930 20156
rect 2930 20100 2986 20156
rect 2986 20100 2990 20156
rect 2926 20096 2990 20100
rect 3006 20156 3070 20160
rect 3006 20100 3010 20156
rect 3010 20100 3066 20156
rect 3066 20100 3070 20156
rect 3006 20096 3070 20100
rect 3086 20156 3150 20160
rect 3086 20100 3090 20156
rect 3090 20100 3146 20156
rect 3146 20100 3150 20156
rect 3086 20096 3150 20100
rect 3166 20156 3230 20160
rect 3166 20100 3170 20156
rect 3170 20100 3226 20156
rect 3226 20100 3230 20156
rect 3166 20096 3230 20100
rect 6874 20156 6938 20160
rect 6874 20100 6878 20156
rect 6878 20100 6934 20156
rect 6934 20100 6938 20156
rect 6874 20096 6938 20100
rect 6954 20156 7018 20160
rect 6954 20100 6958 20156
rect 6958 20100 7014 20156
rect 7014 20100 7018 20156
rect 6954 20096 7018 20100
rect 7034 20156 7098 20160
rect 7034 20100 7038 20156
rect 7038 20100 7094 20156
rect 7094 20100 7098 20156
rect 7034 20096 7098 20100
rect 7114 20156 7178 20160
rect 7114 20100 7118 20156
rect 7118 20100 7174 20156
rect 7174 20100 7178 20156
rect 7114 20096 7178 20100
rect 10822 20156 10886 20160
rect 10822 20100 10826 20156
rect 10826 20100 10882 20156
rect 10882 20100 10886 20156
rect 10822 20096 10886 20100
rect 10902 20156 10966 20160
rect 10902 20100 10906 20156
rect 10906 20100 10962 20156
rect 10962 20100 10966 20156
rect 10902 20096 10966 20100
rect 10982 20156 11046 20160
rect 10982 20100 10986 20156
rect 10986 20100 11042 20156
rect 11042 20100 11046 20156
rect 10982 20096 11046 20100
rect 11062 20156 11126 20160
rect 11062 20100 11066 20156
rect 11066 20100 11122 20156
rect 11122 20100 11126 20156
rect 11062 20096 11126 20100
rect 14770 20156 14834 20160
rect 14770 20100 14774 20156
rect 14774 20100 14830 20156
rect 14830 20100 14834 20156
rect 14770 20096 14834 20100
rect 14850 20156 14914 20160
rect 14850 20100 14854 20156
rect 14854 20100 14910 20156
rect 14910 20100 14914 20156
rect 14850 20096 14914 20100
rect 14930 20156 14994 20160
rect 14930 20100 14934 20156
rect 14934 20100 14990 20156
rect 14990 20100 14994 20156
rect 14930 20096 14994 20100
rect 15010 20156 15074 20160
rect 15010 20100 15014 20156
rect 15014 20100 15070 20156
rect 15070 20100 15074 20156
rect 15010 20096 15074 20100
rect 4900 19612 4964 19616
rect 4900 19556 4904 19612
rect 4904 19556 4960 19612
rect 4960 19556 4964 19612
rect 4900 19552 4964 19556
rect 4980 19612 5044 19616
rect 4980 19556 4984 19612
rect 4984 19556 5040 19612
rect 5040 19556 5044 19612
rect 4980 19552 5044 19556
rect 5060 19612 5124 19616
rect 5060 19556 5064 19612
rect 5064 19556 5120 19612
rect 5120 19556 5124 19612
rect 5060 19552 5124 19556
rect 5140 19612 5204 19616
rect 5140 19556 5144 19612
rect 5144 19556 5200 19612
rect 5200 19556 5204 19612
rect 5140 19552 5204 19556
rect 8848 19612 8912 19616
rect 8848 19556 8852 19612
rect 8852 19556 8908 19612
rect 8908 19556 8912 19612
rect 8848 19552 8912 19556
rect 8928 19612 8992 19616
rect 8928 19556 8932 19612
rect 8932 19556 8988 19612
rect 8988 19556 8992 19612
rect 8928 19552 8992 19556
rect 9008 19612 9072 19616
rect 9008 19556 9012 19612
rect 9012 19556 9068 19612
rect 9068 19556 9072 19612
rect 9008 19552 9072 19556
rect 9088 19612 9152 19616
rect 9088 19556 9092 19612
rect 9092 19556 9148 19612
rect 9148 19556 9152 19612
rect 9088 19552 9152 19556
rect 12796 19612 12860 19616
rect 12796 19556 12800 19612
rect 12800 19556 12856 19612
rect 12856 19556 12860 19612
rect 12796 19552 12860 19556
rect 12876 19612 12940 19616
rect 12876 19556 12880 19612
rect 12880 19556 12936 19612
rect 12936 19556 12940 19612
rect 12876 19552 12940 19556
rect 12956 19612 13020 19616
rect 12956 19556 12960 19612
rect 12960 19556 13016 19612
rect 13016 19556 13020 19612
rect 12956 19552 13020 19556
rect 13036 19612 13100 19616
rect 13036 19556 13040 19612
rect 13040 19556 13096 19612
rect 13096 19556 13100 19612
rect 13036 19552 13100 19556
rect 4476 19212 4540 19276
rect 2926 19068 2990 19072
rect 2926 19012 2930 19068
rect 2930 19012 2986 19068
rect 2986 19012 2990 19068
rect 2926 19008 2990 19012
rect 3006 19068 3070 19072
rect 3006 19012 3010 19068
rect 3010 19012 3066 19068
rect 3066 19012 3070 19068
rect 3006 19008 3070 19012
rect 3086 19068 3150 19072
rect 3086 19012 3090 19068
rect 3090 19012 3146 19068
rect 3146 19012 3150 19068
rect 3086 19008 3150 19012
rect 3166 19068 3230 19072
rect 3166 19012 3170 19068
rect 3170 19012 3226 19068
rect 3226 19012 3230 19068
rect 3166 19008 3230 19012
rect 6874 19068 6938 19072
rect 6874 19012 6878 19068
rect 6878 19012 6934 19068
rect 6934 19012 6938 19068
rect 6874 19008 6938 19012
rect 6954 19068 7018 19072
rect 6954 19012 6958 19068
rect 6958 19012 7014 19068
rect 7014 19012 7018 19068
rect 6954 19008 7018 19012
rect 7034 19068 7098 19072
rect 7034 19012 7038 19068
rect 7038 19012 7094 19068
rect 7094 19012 7098 19068
rect 7034 19008 7098 19012
rect 7114 19068 7178 19072
rect 7114 19012 7118 19068
rect 7118 19012 7174 19068
rect 7174 19012 7178 19068
rect 7114 19008 7178 19012
rect 10822 19068 10886 19072
rect 10822 19012 10826 19068
rect 10826 19012 10882 19068
rect 10882 19012 10886 19068
rect 10822 19008 10886 19012
rect 10902 19068 10966 19072
rect 10902 19012 10906 19068
rect 10906 19012 10962 19068
rect 10962 19012 10966 19068
rect 10902 19008 10966 19012
rect 10982 19068 11046 19072
rect 10982 19012 10986 19068
rect 10986 19012 11042 19068
rect 11042 19012 11046 19068
rect 10982 19008 11046 19012
rect 11062 19068 11126 19072
rect 11062 19012 11066 19068
rect 11066 19012 11122 19068
rect 11122 19012 11126 19068
rect 11062 19008 11126 19012
rect 14770 19068 14834 19072
rect 14770 19012 14774 19068
rect 14774 19012 14830 19068
rect 14830 19012 14834 19068
rect 14770 19008 14834 19012
rect 14850 19068 14914 19072
rect 14850 19012 14854 19068
rect 14854 19012 14910 19068
rect 14910 19012 14914 19068
rect 14850 19008 14914 19012
rect 14930 19068 14994 19072
rect 14930 19012 14934 19068
rect 14934 19012 14990 19068
rect 14990 19012 14994 19068
rect 14930 19008 14994 19012
rect 15010 19068 15074 19072
rect 15010 19012 15014 19068
rect 15014 19012 15070 19068
rect 15070 19012 15074 19068
rect 15010 19008 15074 19012
rect 4660 18804 4724 18868
rect 5764 18668 5828 18732
rect 2452 18532 2516 18596
rect 4900 18524 4964 18528
rect 4900 18468 4904 18524
rect 4904 18468 4960 18524
rect 4960 18468 4964 18524
rect 4900 18464 4964 18468
rect 4980 18524 5044 18528
rect 4980 18468 4984 18524
rect 4984 18468 5040 18524
rect 5040 18468 5044 18524
rect 4980 18464 5044 18468
rect 5060 18524 5124 18528
rect 5060 18468 5064 18524
rect 5064 18468 5120 18524
rect 5120 18468 5124 18524
rect 5060 18464 5124 18468
rect 5140 18524 5204 18528
rect 5140 18468 5144 18524
rect 5144 18468 5200 18524
rect 5200 18468 5204 18524
rect 5140 18464 5204 18468
rect 8848 18524 8912 18528
rect 8848 18468 8852 18524
rect 8852 18468 8908 18524
rect 8908 18468 8912 18524
rect 8848 18464 8912 18468
rect 8928 18524 8992 18528
rect 8928 18468 8932 18524
rect 8932 18468 8988 18524
rect 8988 18468 8992 18524
rect 8928 18464 8992 18468
rect 9008 18524 9072 18528
rect 9008 18468 9012 18524
rect 9012 18468 9068 18524
rect 9068 18468 9072 18524
rect 9008 18464 9072 18468
rect 9088 18524 9152 18528
rect 9088 18468 9092 18524
rect 9092 18468 9148 18524
rect 9148 18468 9152 18524
rect 9088 18464 9152 18468
rect 1716 18260 1780 18324
rect 8708 18396 8772 18460
rect 5948 18260 6012 18324
rect 7788 18260 7852 18324
rect 12796 18524 12860 18528
rect 12796 18468 12800 18524
rect 12800 18468 12856 18524
rect 12856 18468 12860 18524
rect 12796 18464 12860 18468
rect 12876 18524 12940 18528
rect 12876 18468 12880 18524
rect 12880 18468 12936 18524
rect 12936 18468 12940 18524
rect 12876 18464 12940 18468
rect 12956 18524 13020 18528
rect 12956 18468 12960 18524
rect 12960 18468 13016 18524
rect 13016 18468 13020 18524
rect 12956 18464 13020 18468
rect 13036 18524 13100 18528
rect 13036 18468 13040 18524
rect 13040 18468 13096 18524
rect 13096 18468 13100 18524
rect 13036 18464 13100 18468
rect 11468 18396 11532 18460
rect 16804 18260 16868 18324
rect 4108 18048 4172 18052
rect 4108 17992 4122 18048
rect 4122 17992 4172 18048
rect 4108 17988 4172 17992
rect 2926 17980 2990 17984
rect 2926 17924 2930 17980
rect 2930 17924 2986 17980
rect 2986 17924 2990 17980
rect 2926 17920 2990 17924
rect 3006 17980 3070 17984
rect 3006 17924 3010 17980
rect 3010 17924 3066 17980
rect 3066 17924 3070 17980
rect 3006 17920 3070 17924
rect 3086 17980 3150 17984
rect 3086 17924 3090 17980
rect 3090 17924 3146 17980
rect 3146 17924 3150 17980
rect 3086 17920 3150 17924
rect 3166 17980 3230 17984
rect 3166 17924 3170 17980
rect 3170 17924 3226 17980
rect 3226 17924 3230 17980
rect 3166 17920 3230 17924
rect 12572 18124 12636 18188
rect 6132 17988 6196 18052
rect 9260 17988 9324 18052
rect 9812 17988 9876 18052
rect 6874 17980 6938 17984
rect 6874 17924 6878 17980
rect 6878 17924 6934 17980
rect 6934 17924 6938 17980
rect 6874 17920 6938 17924
rect 6954 17980 7018 17984
rect 6954 17924 6958 17980
rect 6958 17924 7014 17980
rect 7014 17924 7018 17980
rect 6954 17920 7018 17924
rect 7034 17980 7098 17984
rect 7034 17924 7038 17980
rect 7038 17924 7094 17980
rect 7094 17924 7098 17980
rect 7034 17920 7098 17924
rect 7114 17980 7178 17984
rect 7114 17924 7118 17980
rect 7118 17924 7174 17980
rect 7174 17924 7178 17980
rect 7114 17920 7178 17924
rect 10822 17980 10886 17984
rect 10822 17924 10826 17980
rect 10826 17924 10882 17980
rect 10882 17924 10886 17980
rect 10822 17920 10886 17924
rect 10902 17980 10966 17984
rect 10902 17924 10906 17980
rect 10906 17924 10962 17980
rect 10962 17924 10966 17980
rect 10902 17920 10966 17924
rect 10982 17980 11046 17984
rect 10982 17924 10986 17980
rect 10986 17924 11042 17980
rect 11042 17924 11046 17980
rect 10982 17920 11046 17924
rect 11062 17980 11126 17984
rect 11062 17924 11066 17980
rect 11066 17924 11122 17980
rect 11122 17924 11126 17980
rect 11062 17920 11126 17924
rect 14770 17980 14834 17984
rect 14770 17924 14774 17980
rect 14774 17924 14830 17980
rect 14830 17924 14834 17980
rect 14770 17920 14834 17924
rect 14850 17980 14914 17984
rect 14850 17924 14854 17980
rect 14854 17924 14910 17980
rect 14910 17924 14914 17980
rect 14850 17920 14914 17924
rect 14930 17980 14994 17984
rect 14930 17924 14934 17980
rect 14934 17924 14990 17980
rect 14990 17924 14994 17980
rect 14930 17920 14994 17924
rect 15010 17980 15074 17984
rect 15010 17924 15014 17980
rect 15014 17924 15070 17980
rect 15070 17924 15074 17980
rect 15010 17920 15074 17924
rect 8156 17852 8220 17916
rect 11652 17444 11716 17508
rect 4900 17436 4964 17440
rect 4900 17380 4904 17436
rect 4904 17380 4960 17436
rect 4960 17380 4964 17436
rect 4900 17376 4964 17380
rect 4980 17436 5044 17440
rect 4980 17380 4984 17436
rect 4984 17380 5040 17436
rect 5040 17380 5044 17436
rect 4980 17376 5044 17380
rect 5060 17436 5124 17440
rect 5060 17380 5064 17436
rect 5064 17380 5120 17436
rect 5120 17380 5124 17436
rect 5060 17376 5124 17380
rect 5140 17436 5204 17440
rect 5140 17380 5144 17436
rect 5144 17380 5200 17436
rect 5200 17380 5204 17436
rect 5140 17376 5204 17380
rect 8848 17436 8912 17440
rect 8848 17380 8852 17436
rect 8852 17380 8908 17436
rect 8908 17380 8912 17436
rect 8848 17376 8912 17380
rect 8928 17436 8992 17440
rect 8928 17380 8932 17436
rect 8932 17380 8988 17436
rect 8988 17380 8992 17436
rect 8928 17376 8992 17380
rect 9008 17436 9072 17440
rect 9008 17380 9012 17436
rect 9012 17380 9068 17436
rect 9068 17380 9072 17436
rect 9008 17376 9072 17380
rect 9088 17436 9152 17440
rect 9088 17380 9092 17436
rect 9092 17380 9148 17436
rect 9148 17380 9152 17436
rect 9088 17376 9152 17380
rect 12796 17436 12860 17440
rect 12796 17380 12800 17436
rect 12800 17380 12856 17436
rect 12856 17380 12860 17436
rect 12796 17376 12860 17380
rect 12876 17436 12940 17440
rect 12876 17380 12880 17436
rect 12880 17380 12936 17436
rect 12936 17380 12940 17436
rect 12876 17376 12940 17380
rect 12956 17436 13020 17440
rect 12956 17380 12960 17436
rect 12960 17380 13016 17436
rect 13016 17380 13020 17436
rect 12956 17376 13020 17380
rect 13036 17436 13100 17440
rect 13036 17380 13040 17436
rect 13040 17380 13096 17436
rect 13096 17380 13100 17436
rect 13036 17376 13100 17380
rect 10548 17308 10612 17372
rect 3924 17172 3988 17236
rect 6500 17036 6564 17100
rect 9444 17036 9508 17100
rect 9812 17036 9876 17100
rect 14044 17036 14108 17100
rect 7972 16900 8036 16964
rect 2926 16892 2990 16896
rect 2926 16836 2930 16892
rect 2930 16836 2986 16892
rect 2986 16836 2990 16892
rect 2926 16832 2990 16836
rect 3006 16892 3070 16896
rect 3006 16836 3010 16892
rect 3010 16836 3066 16892
rect 3066 16836 3070 16892
rect 3006 16832 3070 16836
rect 3086 16892 3150 16896
rect 3086 16836 3090 16892
rect 3090 16836 3146 16892
rect 3146 16836 3150 16892
rect 3086 16832 3150 16836
rect 3166 16892 3230 16896
rect 3166 16836 3170 16892
rect 3170 16836 3226 16892
rect 3226 16836 3230 16892
rect 3166 16832 3230 16836
rect 6874 16892 6938 16896
rect 6874 16836 6878 16892
rect 6878 16836 6934 16892
rect 6934 16836 6938 16892
rect 6874 16832 6938 16836
rect 6954 16892 7018 16896
rect 6954 16836 6958 16892
rect 6958 16836 7014 16892
rect 7014 16836 7018 16892
rect 6954 16832 7018 16836
rect 7034 16892 7098 16896
rect 7034 16836 7038 16892
rect 7038 16836 7094 16892
rect 7094 16836 7098 16892
rect 7034 16832 7098 16836
rect 7114 16892 7178 16896
rect 7114 16836 7118 16892
rect 7118 16836 7174 16892
rect 7174 16836 7178 16892
rect 7114 16832 7178 16836
rect 10822 16892 10886 16896
rect 10822 16836 10826 16892
rect 10826 16836 10882 16892
rect 10882 16836 10886 16892
rect 10822 16832 10886 16836
rect 10902 16892 10966 16896
rect 10902 16836 10906 16892
rect 10906 16836 10962 16892
rect 10962 16836 10966 16892
rect 10902 16832 10966 16836
rect 10982 16892 11046 16896
rect 10982 16836 10986 16892
rect 10986 16836 11042 16892
rect 11042 16836 11046 16892
rect 10982 16832 11046 16836
rect 11062 16892 11126 16896
rect 11062 16836 11066 16892
rect 11066 16836 11122 16892
rect 11122 16836 11126 16892
rect 11062 16832 11126 16836
rect 14770 16892 14834 16896
rect 14770 16836 14774 16892
rect 14774 16836 14830 16892
rect 14830 16836 14834 16892
rect 14770 16832 14834 16836
rect 14850 16892 14914 16896
rect 14850 16836 14854 16892
rect 14854 16836 14910 16892
rect 14910 16836 14914 16892
rect 14850 16832 14914 16836
rect 14930 16892 14994 16896
rect 14930 16836 14934 16892
rect 14934 16836 14990 16892
rect 14990 16836 14994 16892
rect 14930 16832 14994 16836
rect 15010 16892 15074 16896
rect 15010 16836 15014 16892
rect 15014 16836 15070 16892
rect 15070 16836 15074 16892
rect 15010 16832 15074 16836
rect 5396 16824 5460 16828
rect 5396 16768 5446 16824
rect 5446 16768 5460 16824
rect 5396 16764 5460 16768
rect 8708 16764 8772 16828
rect 2452 16628 2516 16692
rect 7604 16628 7668 16692
rect 8524 16628 8588 16692
rect 2268 16492 2332 16556
rect 3372 16492 3436 16556
rect 5580 16492 5644 16556
rect 7420 16552 7484 16556
rect 7420 16496 7434 16552
rect 7434 16496 7484 16552
rect 7420 16492 7484 16496
rect 2636 16356 2700 16420
rect 6684 16416 6748 16420
rect 6684 16360 6734 16416
rect 6734 16360 6748 16416
rect 6684 16356 6748 16360
rect 4900 16348 4964 16352
rect 4900 16292 4904 16348
rect 4904 16292 4960 16348
rect 4960 16292 4964 16348
rect 4900 16288 4964 16292
rect 4980 16348 5044 16352
rect 4980 16292 4984 16348
rect 4984 16292 5040 16348
rect 5040 16292 5044 16348
rect 4980 16288 5044 16292
rect 5060 16348 5124 16352
rect 5060 16292 5064 16348
rect 5064 16292 5120 16348
rect 5120 16292 5124 16348
rect 5060 16288 5124 16292
rect 5140 16348 5204 16352
rect 5140 16292 5144 16348
rect 5144 16292 5200 16348
rect 5200 16292 5204 16348
rect 5140 16288 5204 16292
rect 6316 16220 6380 16284
rect 9812 16356 9876 16420
rect 9996 16416 10060 16420
rect 9996 16360 10010 16416
rect 10010 16360 10060 16416
rect 9996 16356 10060 16360
rect 12020 16356 12084 16420
rect 8848 16348 8912 16352
rect 8848 16292 8852 16348
rect 8852 16292 8908 16348
rect 8908 16292 8912 16348
rect 8848 16288 8912 16292
rect 8928 16348 8992 16352
rect 8928 16292 8932 16348
rect 8932 16292 8988 16348
rect 8988 16292 8992 16348
rect 8928 16288 8992 16292
rect 9008 16348 9072 16352
rect 9008 16292 9012 16348
rect 9012 16292 9068 16348
rect 9068 16292 9072 16348
rect 9008 16288 9072 16292
rect 9088 16348 9152 16352
rect 9088 16292 9092 16348
rect 9092 16292 9148 16348
rect 9148 16292 9152 16348
rect 9088 16288 9152 16292
rect 12796 16348 12860 16352
rect 12796 16292 12800 16348
rect 12800 16292 12856 16348
rect 12856 16292 12860 16348
rect 12796 16288 12860 16292
rect 12876 16348 12940 16352
rect 12876 16292 12880 16348
rect 12880 16292 12936 16348
rect 12936 16292 12940 16348
rect 12876 16288 12940 16292
rect 12956 16348 13020 16352
rect 12956 16292 12960 16348
rect 12960 16292 13016 16348
rect 13016 16292 13020 16348
rect 12956 16288 13020 16292
rect 13036 16348 13100 16352
rect 13036 16292 13040 16348
rect 13040 16292 13096 16348
rect 13096 16292 13100 16348
rect 13036 16288 13100 16292
rect 2452 15948 2516 16012
rect 11836 15948 11900 16012
rect 4292 15812 4356 15876
rect 5396 15812 5460 15876
rect 8708 15812 8772 15876
rect 2926 15804 2990 15808
rect 2926 15748 2930 15804
rect 2930 15748 2986 15804
rect 2986 15748 2990 15804
rect 2926 15744 2990 15748
rect 3006 15804 3070 15808
rect 3006 15748 3010 15804
rect 3010 15748 3066 15804
rect 3066 15748 3070 15804
rect 3006 15744 3070 15748
rect 3086 15804 3150 15808
rect 3086 15748 3090 15804
rect 3090 15748 3146 15804
rect 3146 15748 3150 15804
rect 3086 15744 3150 15748
rect 3166 15804 3230 15808
rect 3166 15748 3170 15804
rect 3170 15748 3226 15804
rect 3226 15748 3230 15804
rect 3166 15744 3230 15748
rect 6874 15804 6938 15808
rect 6874 15748 6878 15804
rect 6878 15748 6934 15804
rect 6934 15748 6938 15804
rect 6874 15744 6938 15748
rect 6954 15804 7018 15808
rect 6954 15748 6958 15804
rect 6958 15748 7014 15804
rect 7014 15748 7018 15804
rect 6954 15744 7018 15748
rect 7034 15804 7098 15808
rect 7034 15748 7038 15804
rect 7038 15748 7094 15804
rect 7094 15748 7098 15804
rect 7034 15744 7098 15748
rect 7114 15804 7178 15808
rect 7114 15748 7118 15804
rect 7118 15748 7174 15804
rect 7174 15748 7178 15804
rect 7114 15744 7178 15748
rect 10822 15804 10886 15808
rect 10822 15748 10826 15804
rect 10826 15748 10882 15804
rect 10882 15748 10886 15804
rect 10822 15744 10886 15748
rect 10902 15804 10966 15808
rect 10902 15748 10906 15804
rect 10906 15748 10962 15804
rect 10962 15748 10966 15804
rect 10902 15744 10966 15748
rect 10982 15804 11046 15808
rect 10982 15748 10986 15804
rect 10986 15748 11042 15804
rect 11042 15748 11046 15804
rect 10982 15744 11046 15748
rect 11062 15804 11126 15808
rect 11062 15748 11066 15804
rect 11066 15748 11122 15804
rect 11122 15748 11126 15804
rect 11062 15744 11126 15748
rect 14770 15804 14834 15808
rect 14770 15748 14774 15804
rect 14774 15748 14830 15804
rect 14830 15748 14834 15804
rect 14770 15744 14834 15748
rect 14850 15804 14914 15808
rect 14850 15748 14854 15804
rect 14854 15748 14910 15804
rect 14910 15748 14914 15804
rect 14850 15744 14914 15748
rect 14930 15804 14994 15808
rect 14930 15748 14934 15804
rect 14934 15748 14990 15804
rect 14990 15748 14994 15804
rect 14930 15744 14994 15748
rect 15010 15804 15074 15808
rect 15010 15748 15014 15804
rect 15014 15748 15070 15804
rect 15070 15748 15074 15804
rect 15010 15744 15074 15748
rect 7282 15676 7346 15740
rect 7972 15676 8036 15740
rect 3556 15540 3620 15604
rect 8340 15540 8404 15604
rect 15884 15540 15948 15604
rect 9812 15404 9876 15468
rect 13860 15404 13924 15468
rect 1900 15268 1964 15332
rect 5396 15268 5460 15332
rect 7604 15268 7668 15332
rect 4900 15260 4964 15264
rect 4900 15204 4904 15260
rect 4904 15204 4960 15260
rect 4960 15204 4964 15260
rect 4900 15200 4964 15204
rect 4980 15260 5044 15264
rect 4980 15204 4984 15260
rect 4984 15204 5040 15260
rect 5040 15204 5044 15260
rect 4980 15200 5044 15204
rect 5060 15260 5124 15264
rect 5060 15204 5064 15260
rect 5064 15204 5120 15260
rect 5120 15204 5124 15260
rect 5060 15200 5124 15204
rect 5140 15260 5204 15264
rect 5140 15204 5144 15260
rect 5144 15204 5200 15260
rect 5200 15204 5204 15260
rect 5140 15200 5204 15204
rect 6132 15192 6196 15196
rect 6132 15136 6146 15192
rect 6146 15136 6196 15192
rect 6132 15132 6196 15136
rect 6132 14996 6196 15060
rect 8848 15260 8912 15264
rect 8848 15204 8852 15260
rect 8852 15204 8908 15260
rect 8908 15204 8912 15260
rect 8848 15200 8912 15204
rect 8928 15260 8992 15264
rect 8928 15204 8932 15260
rect 8932 15204 8988 15260
rect 8988 15204 8992 15260
rect 8928 15200 8992 15204
rect 9008 15260 9072 15264
rect 9008 15204 9012 15260
rect 9012 15204 9068 15260
rect 9068 15204 9072 15260
rect 9008 15200 9072 15204
rect 9088 15260 9152 15264
rect 9088 15204 9092 15260
rect 9092 15204 9148 15260
rect 9148 15204 9152 15260
rect 9088 15200 9152 15204
rect 12796 15260 12860 15264
rect 12796 15204 12800 15260
rect 12800 15204 12856 15260
rect 12856 15204 12860 15260
rect 12796 15200 12860 15204
rect 12876 15260 12940 15264
rect 12876 15204 12880 15260
rect 12880 15204 12936 15260
rect 12936 15204 12940 15260
rect 12876 15200 12940 15204
rect 12956 15260 13020 15264
rect 12956 15204 12960 15260
rect 12960 15204 13016 15260
rect 13016 15204 13020 15260
rect 12956 15200 13020 15204
rect 13036 15260 13100 15264
rect 13036 15204 13040 15260
rect 13040 15204 13096 15260
rect 13096 15204 13100 15260
rect 13036 15200 13100 15204
rect 11284 15132 11348 15196
rect 12388 15132 12452 15196
rect 9812 14996 9876 15060
rect 10180 14996 10244 15060
rect 15516 14996 15580 15060
rect 2926 14716 2990 14720
rect 2926 14660 2930 14716
rect 2930 14660 2986 14716
rect 2986 14660 2990 14716
rect 2926 14656 2990 14660
rect 3006 14716 3070 14720
rect 3006 14660 3010 14716
rect 3010 14660 3066 14716
rect 3066 14660 3070 14716
rect 3006 14656 3070 14660
rect 3086 14716 3150 14720
rect 3086 14660 3090 14716
rect 3090 14660 3146 14716
rect 3146 14660 3150 14716
rect 3086 14656 3150 14660
rect 3166 14716 3230 14720
rect 3166 14660 3170 14716
rect 3170 14660 3226 14716
rect 3226 14660 3230 14716
rect 3166 14656 3230 14660
rect 2268 14588 2332 14652
rect 3740 14860 3804 14924
rect 4476 14860 4540 14924
rect 3740 14724 3804 14788
rect 6874 14716 6938 14720
rect 6874 14660 6878 14716
rect 6878 14660 6934 14716
rect 6934 14660 6938 14716
rect 6874 14656 6938 14660
rect 6954 14716 7018 14720
rect 6954 14660 6958 14716
rect 6958 14660 7014 14716
rect 7014 14660 7018 14716
rect 6954 14656 7018 14660
rect 7034 14716 7098 14720
rect 7034 14660 7038 14716
rect 7038 14660 7094 14716
rect 7094 14660 7098 14716
rect 7034 14656 7098 14660
rect 7114 14716 7178 14720
rect 7114 14660 7118 14716
rect 7118 14660 7174 14716
rect 7174 14660 7178 14716
rect 7114 14656 7178 14660
rect 4476 14648 4540 14652
rect 4476 14592 4526 14648
rect 4526 14592 4540 14648
rect 2268 14316 2332 14380
rect 3556 14316 3620 14380
rect 3556 14180 3620 14244
rect 4476 14588 4540 14592
rect 7972 14724 8036 14788
rect 9260 14724 9324 14788
rect 16436 14860 16500 14924
rect 13676 14724 13740 14788
rect 10822 14716 10886 14720
rect 10822 14660 10826 14716
rect 10826 14660 10882 14716
rect 10882 14660 10886 14716
rect 10822 14656 10886 14660
rect 10902 14716 10966 14720
rect 10902 14660 10906 14716
rect 10906 14660 10962 14716
rect 10962 14660 10966 14716
rect 10902 14656 10966 14660
rect 10982 14716 11046 14720
rect 10982 14660 10986 14716
rect 10986 14660 11042 14716
rect 11042 14660 11046 14716
rect 10982 14656 11046 14660
rect 11062 14716 11126 14720
rect 11062 14660 11066 14716
rect 11066 14660 11122 14716
rect 11122 14660 11126 14716
rect 11062 14656 11126 14660
rect 14770 14716 14834 14720
rect 14770 14660 14774 14716
rect 14774 14660 14830 14716
rect 14830 14660 14834 14716
rect 14770 14656 14834 14660
rect 14850 14716 14914 14720
rect 14850 14660 14854 14716
rect 14854 14660 14910 14716
rect 14910 14660 14914 14716
rect 14850 14656 14914 14660
rect 14930 14716 14994 14720
rect 14930 14660 14934 14716
rect 14934 14660 14990 14716
rect 14990 14660 14994 14716
rect 14930 14656 14994 14660
rect 15010 14716 15074 14720
rect 15010 14660 15014 14716
rect 15014 14660 15070 14716
rect 15070 14660 15074 14716
rect 15010 14656 15074 14660
rect 12204 14588 12268 14652
rect 3924 14316 3988 14380
rect 13492 14512 13556 14516
rect 13492 14456 13542 14512
rect 13542 14456 13556 14512
rect 13492 14452 13556 14456
rect 4900 14172 4964 14176
rect 4900 14116 4904 14172
rect 4904 14116 4960 14172
rect 4960 14116 4964 14172
rect 4900 14112 4964 14116
rect 4980 14172 5044 14176
rect 4980 14116 4984 14172
rect 4984 14116 5040 14172
rect 5040 14116 5044 14172
rect 4980 14112 5044 14116
rect 5060 14172 5124 14176
rect 5060 14116 5064 14172
rect 5064 14116 5120 14172
rect 5120 14116 5124 14172
rect 5060 14112 5124 14116
rect 5140 14172 5204 14176
rect 5140 14116 5144 14172
rect 5144 14116 5200 14172
rect 5200 14116 5204 14172
rect 5140 14112 5204 14116
rect 2926 13628 2990 13632
rect 2926 13572 2930 13628
rect 2930 13572 2986 13628
rect 2986 13572 2990 13628
rect 2926 13568 2990 13572
rect 3006 13628 3070 13632
rect 3006 13572 3010 13628
rect 3010 13572 3066 13628
rect 3066 13572 3070 13628
rect 3006 13568 3070 13572
rect 3086 13628 3150 13632
rect 3086 13572 3090 13628
rect 3090 13572 3146 13628
rect 3146 13572 3150 13628
rect 3086 13568 3150 13572
rect 3166 13628 3230 13632
rect 3166 13572 3170 13628
rect 3170 13572 3226 13628
rect 3226 13572 3230 13628
rect 3166 13568 3230 13572
rect 5948 14044 6012 14108
rect 8848 14172 8912 14176
rect 8848 14116 8852 14172
rect 8852 14116 8908 14172
rect 8908 14116 8912 14172
rect 8848 14112 8912 14116
rect 8928 14172 8992 14176
rect 8928 14116 8932 14172
rect 8932 14116 8988 14172
rect 8988 14116 8992 14172
rect 8928 14112 8992 14116
rect 9008 14172 9072 14176
rect 9008 14116 9012 14172
rect 9012 14116 9068 14172
rect 9068 14116 9072 14172
rect 9008 14112 9072 14116
rect 9088 14172 9152 14176
rect 9088 14116 9092 14172
rect 9092 14116 9148 14172
rect 9148 14116 9152 14172
rect 9088 14112 9152 14116
rect 9628 14316 9692 14380
rect 10364 14180 10428 14244
rect 11284 14180 11348 14244
rect 13308 14180 13372 14244
rect 12796 14172 12860 14176
rect 12796 14116 12800 14172
rect 12800 14116 12856 14172
rect 12856 14116 12860 14172
rect 12796 14112 12860 14116
rect 12876 14172 12940 14176
rect 12876 14116 12880 14172
rect 12880 14116 12936 14172
rect 12936 14116 12940 14172
rect 12876 14112 12940 14116
rect 12956 14172 13020 14176
rect 12956 14116 12960 14172
rect 12960 14116 13016 14172
rect 13016 14116 13020 14172
rect 12956 14112 13020 14116
rect 13036 14172 13100 14176
rect 13036 14116 13040 14172
rect 13040 14116 13096 14172
rect 13096 14116 13100 14172
rect 13036 14112 13100 14116
rect 14412 13908 14476 13972
rect 8708 13772 8772 13836
rect 4476 13636 4540 13700
rect 5580 13696 5644 13700
rect 5580 13640 5630 13696
rect 5630 13640 5644 13696
rect 5580 13636 5644 13640
rect 6874 13628 6938 13632
rect 6874 13572 6878 13628
rect 6878 13572 6934 13628
rect 6934 13572 6938 13628
rect 6874 13568 6938 13572
rect 6954 13628 7018 13632
rect 6954 13572 6958 13628
rect 6958 13572 7014 13628
rect 7014 13572 7018 13628
rect 6954 13568 7018 13572
rect 7034 13628 7098 13632
rect 7034 13572 7038 13628
rect 7038 13572 7094 13628
rect 7094 13572 7098 13628
rect 7034 13568 7098 13572
rect 7114 13628 7178 13632
rect 7114 13572 7118 13628
rect 7118 13572 7174 13628
rect 7174 13572 7178 13628
rect 7114 13568 7178 13572
rect 5580 13500 5644 13564
rect 7788 13500 7852 13564
rect 4476 13424 4540 13428
rect 4476 13368 4526 13424
rect 4526 13368 4540 13424
rect 4476 13364 4540 13368
rect 11284 13636 11348 13700
rect 14596 13636 14660 13700
rect 10822 13628 10886 13632
rect 10822 13572 10826 13628
rect 10826 13572 10882 13628
rect 10882 13572 10886 13628
rect 10822 13568 10886 13572
rect 10902 13628 10966 13632
rect 10902 13572 10906 13628
rect 10906 13572 10962 13628
rect 10962 13572 10966 13628
rect 10902 13568 10966 13572
rect 10982 13628 11046 13632
rect 10982 13572 10986 13628
rect 10986 13572 11042 13628
rect 11042 13572 11046 13628
rect 10982 13568 11046 13572
rect 11062 13628 11126 13632
rect 11062 13572 11066 13628
rect 11066 13572 11122 13628
rect 11122 13572 11126 13628
rect 11062 13568 11126 13572
rect 14770 13628 14834 13632
rect 14770 13572 14774 13628
rect 14774 13572 14830 13628
rect 14830 13572 14834 13628
rect 14770 13568 14834 13572
rect 14850 13628 14914 13632
rect 14850 13572 14854 13628
rect 14854 13572 14910 13628
rect 14910 13572 14914 13628
rect 14850 13568 14914 13572
rect 14930 13628 14994 13632
rect 14930 13572 14934 13628
rect 14934 13572 14990 13628
rect 14990 13572 14994 13628
rect 14930 13568 14994 13572
rect 15010 13628 15074 13632
rect 15010 13572 15014 13628
rect 15014 13572 15070 13628
rect 15070 13572 15074 13628
rect 15010 13568 15074 13572
rect 8708 13500 8772 13564
rect 13170 13500 13234 13564
rect 14228 13500 14292 13564
rect 15332 13560 15396 13564
rect 15332 13504 15382 13560
rect 15382 13504 15396 13560
rect 15332 13500 15396 13504
rect 15148 13228 15212 13292
rect 15700 13288 15764 13292
rect 15700 13232 15714 13288
rect 15714 13232 15764 13288
rect 15700 13228 15764 13232
rect 5948 13092 6012 13156
rect 4900 13084 4964 13088
rect 4900 13028 4904 13084
rect 4904 13028 4960 13084
rect 4960 13028 4964 13084
rect 4900 13024 4964 13028
rect 4980 13084 5044 13088
rect 4980 13028 4984 13084
rect 4984 13028 5040 13084
rect 5040 13028 5044 13084
rect 4980 13024 5044 13028
rect 5060 13084 5124 13088
rect 5060 13028 5064 13084
rect 5064 13028 5120 13084
rect 5120 13028 5124 13084
rect 5060 13024 5124 13028
rect 5140 13084 5204 13088
rect 5140 13028 5144 13084
rect 5144 13028 5200 13084
rect 5200 13028 5204 13084
rect 5140 13024 5204 13028
rect 11652 13092 11716 13156
rect 8848 13084 8912 13088
rect 8848 13028 8852 13084
rect 8852 13028 8908 13084
rect 8908 13028 8912 13084
rect 8848 13024 8912 13028
rect 8928 13084 8992 13088
rect 8928 13028 8932 13084
rect 8932 13028 8988 13084
rect 8988 13028 8992 13084
rect 8928 13024 8992 13028
rect 9008 13084 9072 13088
rect 9008 13028 9012 13084
rect 9012 13028 9068 13084
rect 9068 13028 9072 13084
rect 9008 13024 9072 13028
rect 9088 13084 9152 13088
rect 9088 13028 9092 13084
rect 9092 13028 9148 13084
rect 9148 13028 9152 13084
rect 9088 13024 9152 13028
rect 3740 12956 3804 13020
rect 4660 13016 4724 13020
rect 4660 12960 4710 13016
rect 4710 12960 4724 13016
rect 4660 12956 4724 12960
rect 3556 12820 3620 12884
rect 3924 12820 3988 12884
rect 6132 12820 6196 12884
rect 4660 12684 4724 12748
rect 5764 12684 5828 12748
rect 8156 12956 8220 13020
rect 11652 12956 11716 13020
rect 12796 13084 12860 13088
rect 12796 13028 12800 13084
rect 12800 13028 12856 13084
rect 12856 13028 12860 13084
rect 12796 13024 12860 13028
rect 12876 13084 12940 13088
rect 12876 13028 12880 13084
rect 12880 13028 12936 13084
rect 12936 13028 12940 13084
rect 12876 13024 12940 13028
rect 12956 13084 13020 13088
rect 12956 13028 12960 13084
rect 12960 13028 13016 13084
rect 13016 13028 13020 13084
rect 12956 13024 13020 13028
rect 13036 13084 13100 13088
rect 13036 13028 13040 13084
rect 13040 13028 13096 13084
rect 13096 13028 13100 13084
rect 13036 13024 13100 13028
rect 16068 12956 16132 13020
rect 3556 12608 3620 12612
rect 3556 12552 3606 12608
rect 3606 12552 3620 12608
rect 3556 12548 3620 12552
rect 3740 12548 3804 12612
rect 9444 12684 9508 12748
rect 7788 12548 7852 12612
rect 8156 12548 8220 12612
rect 9444 12548 9508 12612
rect 2926 12540 2990 12544
rect 2926 12484 2930 12540
rect 2930 12484 2986 12540
rect 2986 12484 2990 12540
rect 2926 12480 2990 12484
rect 3006 12540 3070 12544
rect 3006 12484 3010 12540
rect 3010 12484 3066 12540
rect 3066 12484 3070 12540
rect 3006 12480 3070 12484
rect 3086 12540 3150 12544
rect 3086 12484 3090 12540
rect 3090 12484 3146 12540
rect 3146 12484 3150 12540
rect 3086 12480 3150 12484
rect 3166 12540 3230 12544
rect 3166 12484 3170 12540
rect 3170 12484 3226 12540
rect 3226 12484 3230 12540
rect 3166 12480 3230 12484
rect 6874 12540 6938 12544
rect 6874 12484 6878 12540
rect 6878 12484 6934 12540
rect 6934 12484 6938 12540
rect 6874 12480 6938 12484
rect 6954 12540 7018 12544
rect 6954 12484 6958 12540
rect 6958 12484 7014 12540
rect 7014 12484 7018 12540
rect 6954 12480 7018 12484
rect 7034 12540 7098 12544
rect 7034 12484 7038 12540
rect 7038 12484 7094 12540
rect 7094 12484 7098 12540
rect 7034 12480 7098 12484
rect 7114 12540 7178 12544
rect 7114 12484 7118 12540
rect 7118 12484 7174 12540
rect 7174 12484 7178 12540
rect 7114 12480 7178 12484
rect 4292 12412 4356 12476
rect 6500 12412 6564 12476
rect 4292 12276 4356 12340
rect 1716 12140 1780 12204
rect 3740 12140 3804 12204
rect 3740 12004 3804 12068
rect 4292 12004 4356 12068
rect 6684 12200 6748 12204
rect 6684 12144 6734 12200
rect 6734 12144 6748 12200
rect 6684 12140 6748 12144
rect 8708 12412 8772 12476
rect 14044 12820 14108 12884
rect 15516 12880 15580 12884
rect 15516 12824 15530 12880
rect 15530 12824 15580 12880
rect 15516 12820 15580 12824
rect 10822 12540 10886 12544
rect 10822 12484 10826 12540
rect 10826 12484 10882 12540
rect 10882 12484 10886 12540
rect 10822 12480 10886 12484
rect 10902 12540 10966 12544
rect 10902 12484 10906 12540
rect 10906 12484 10962 12540
rect 10962 12484 10966 12540
rect 10902 12480 10966 12484
rect 10982 12540 11046 12544
rect 10982 12484 10986 12540
rect 10986 12484 11042 12540
rect 11042 12484 11046 12540
rect 10982 12480 11046 12484
rect 11062 12540 11126 12544
rect 11062 12484 11066 12540
rect 11066 12484 11122 12540
rect 11122 12484 11126 12540
rect 11062 12480 11126 12484
rect 11468 12412 11532 12476
rect 15516 12548 15580 12612
rect 14770 12540 14834 12544
rect 14770 12484 14774 12540
rect 14774 12484 14830 12540
rect 14830 12484 14834 12540
rect 14770 12480 14834 12484
rect 14850 12540 14914 12544
rect 14850 12484 14854 12540
rect 14854 12484 14910 12540
rect 14910 12484 14914 12540
rect 14850 12480 14914 12484
rect 14930 12540 14994 12544
rect 14930 12484 14934 12540
rect 14934 12484 14990 12540
rect 14990 12484 14994 12540
rect 14930 12480 14994 12484
rect 15010 12540 15074 12544
rect 15010 12484 15014 12540
rect 15014 12484 15070 12540
rect 15070 12484 15074 12540
rect 15010 12480 15074 12484
rect 10364 12276 10428 12340
rect 7972 12140 8036 12204
rect 9812 12200 9876 12204
rect 11468 12276 11532 12340
rect 9812 12144 9826 12200
rect 9826 12144 9876 12200
rect 9812 12140 9876 12144
rect 2636 11928 2700 11932
rect 2636 11872 2650 11928
rect 2650 11872 2700 11928
rect 2636 11868 2700 11872
rect 4292 11868 4356 11932
rect 2268 11792 2332 11796
rect 8708 12004 8772 12068
rect 9812 12004 9876 12068
rect 10364 12004 10428 12068
rect 14044 12140 14108 12204
rect 15148 12140 15212 12204
rect 16252 12140 16316 12204
rect 12388 12004 12452 12068
rect 4900 11996 4964 12000
rect 4900 11940 4904 11996
rect 4904 11940 4960 11996
rect 4960 11940 4964 11996
rect 4900 11936 4964 11940
rect 4980 11996 5044 12000
rect 4980 11940 4984 11996
rect 4984 11940 5040 11996
rect 5040 11940 5044 11996
rect 4980 11936 5044 11940
rect 5060 11996 5124 12000
rect 5060 11940 5064 11996
rect 5064 11940 5120 11996
rect 5120 11940 5124 11996
rect 5060 11936 5124 11940
rect 5140 11996 5204 12000
rect 5140 11940 5144 11996
rect 5144 11940 5200 11996
rect 5200 11940 5204 11996
rect 5140 11936 5204 11940
rect 8848 11996 8912 12000
rect 8848 11940 8852 11996
rect 8852 11940 8908 11996
rect 8908 11940 8912 11996
rect 8848 11936 8912 11940
rect 8928 11996 8992 12000
rect 8928 11940 8932 11996
rect 8932 11940 8988 11996
rect 8988 11940 8992 11996
rect 8928 11936 8992 11940
rect 9008 11996 9072 12000
rect 9008 11940 9012 11996
rect 9012 11940 9068 11996
rect 9068 11940 9072 11996
rect 9008 11936 9072 11940
rect 9088 11996 9152 12000
rect 9088 11940 9092 11996
rect 9092 11940 9148 11996
rect 9148 11940 9152 11996
rect 9088 11936 9152 11940
rect 12796 11996 12860 12000
rect 12796 11940 12800 11996
rect 12800 11940 12856 11996
rect 12856 11940 12860 11996
rect 12796 11936 12860 11940
rect 12876 11996 12940 12000
rect 12876 11940 12880 11996
rect 12880 11940 12936 11996
rect 12936 11940 12940 11996
rect 12876 11936 12940 11940
rect 12956 11996 13020 12000
rect 12956 11940 12960 11996
rect 12960 11940 13016 11996
rect 13016 11940 13020 11996
rect 12956 11936 13020 11940
rect 13036 11996 13100 12000
rect 13036 11940 13040 11996
rect 13040 11940 13096 11996
rect 13096 11940 13100 11996
rect 13036 11936 13100 11940
rect 7282 11868 7346 11932
rect 2268 11736 2282 11792
rect 2282 11736 2332 11792
rect 2268 11732 2332 11736
rect 5396 11732 5460 11796
rect 12388 11928 12452 11932
rect 12388 11872 12402 11928
rect 12402 11872 12452 11928
rect 12388 11868 12452 11872
rect 14044 12004 14108 12068
rect 13860 11732 13924 11796
rect 15148 11732 15212 11796
rect 8524 11596 8588 11660
rect 8708 11596 8772 11660
rect 13860 11596 13924 11660
rect 6316 11460 6380 11524
rect 8156 11460 8220 11524
rect 8524 11460 8588 11524
rect 11836 11460 11900 11524
rect 2926 11452 2990 11456
rect 2926 11396 2930 11452
rect 2930 11396 2986 11452
rect 2986 11396 2990 11452
rect 2926 11392 2990 11396
rect 3006 11452 3070 11456
rect 3006 11396 3010 11452
rect 3010 11396 3066 11452
rect 3066 11396 3070 11452
rect 3006 11392 3070 11396
rect 3086 11452 3150 11456
rect 3086 11396 3090 11452
rect 3090 11396 3146 11452
rect 3146 11396 3150 11452
rect 3086 11392 3150 11396
rect 3166 11452 3230 11456
rect 3166 11396 3170 11452
rect 3170 11396 3226 11452
rect 3226 11396 3230 11452
rect 3166 11392 3230 11396
rect 6874 11452 6938 11456
rect 6874 11396 6878 11452
rect 6878 11396 6934 11452
rect 6934 11396 6938 11452
rect 6874 11392 6938 11396
rect 6954 11452 7018 11456
rect 6954 11396 6958 11452
rect 6958 11396 7014 11452
rect 7014 11396 7018 11452
rect 6954 11392 7018 11396
rect 7034 11452 7098 11456
rect 7034 11396 7038 11452
rect 7038 11396 7094 11452
rect 7094 11396 7098 11452
rect 7034 11392 7098 11396
rect 7114 11452 7178 11456
rect 7114 11396 7118 11452
rect 7118 11396 7174 11452
rect 7174 11396 7178 11452
rect 7114 11392 7178 11396
rect 10822 11452 10886 11456
rect 10822 11396 10826 11452
rect 10826 11396 10882 11452
rect 10882 11396 10886 11452
rect 10822 11392 10886 11396
rect 10902 11452 10966 11456
rect 10902 11396 10906 11452
rect 10906 11396 10962 11452
rect 10962 11396 10966 11452
rect 10902 11392 10966 11396
rect 10982 11452 11046 11456
rect 10982 11396 10986 11452
rect 10986 11396 11042 11452
rect 11042 11396 11046 11452
rect 10982 11392 11046 11396
rect 11062 11452 11126 11456
rect 11062 11396 11066 11452
rect 11066 11396 11122 11452
rect 11122 11396 11126 11452
rect 11062 11392 11126 11396
rect 13170 11460 13234 11524
rect 14044 11460 14108 11524
rect 3372 11324 3436 11388
rect 3556 11188 3620 11252
rect 4660 11324 4724 11388
rect 9260 11324 9324 11388
rect 15700 11596 15764 11660
rect 14770 11452 14834 11456
rect 14770 11396 14774 11452
rect 14774 11396 14830 11452
rect 14830 11396 14834 11452
rect 14770 11392 14834 11396
rect 14850 11452 14914 11456
rect 14850 11396 14854 11452
rect 14854 11396 14910 11452
rect 14910 11396 14914 11452
rect 14850 11392 14914 11396
rect 14930 11452 14994 11456
rect 14930 11396 14934 11452
rect 14934 11396 14990 11452
rect 14990 11396 14994 11452
rect 14930 11392 14994 11396
rect 15010 11452 15074 11456
rect 15010 11396 15014 11452
rect 15014 11396 15070 11452
rect 15070 11396 15074 11452
rect 15010 11392 15074 11396
rect 5948 11188 6012 11252
rect 8156 11188 8220 11252
rect 2452 11052 2516 11116
rect 11468 11052 11532 11116
rect 3924 10976 3988 10980
rect 3924 10920 3938 10976
rect 3938 10920 3988 10976
rect 3924 10916 3988 10920
rect 4660 10976 4724 10980
rect 4660 10920 4710 10976
rect 4710 10920 4724 10976
rect 4660 10916 4724 10920
rect 8708 10916 8772 10980
rect 10180 10916 10244 10980
rect 11468 10916 11532 10980
rect 4900 10908 4964 10912
rect 4900 10852 4904 10908
rect 4904 10852 4960 10908
rect 4960 10852 4964 10908
rect 4900 10848 4964 10852
rect 4980 10908 5044 10912
rect 4980 10852 4984 10908
rect 4984 10852 5040 10908
rect 5040 10852 5044 10908
rect 4980 10848 5044 10852
rect 5060 10908 5124 10912
rect 5060 10852 5064 10908
rect 5064 10852 5120 10908
rect 5120 10852 5124 10908
rect 5060 10848 5124 10852
rect 5140 10908 5204 10912
rect 5140 10852 5144 10908
rect 5144 10852 5200 10908
rect 5200 10852 5204 10908
rect 5140 10848 5204 10852
rect 8848 10908 8912 10912
rect 8848 10852 8852 10908
rect 8852 10852 8908 10908
rect 8908 10852 8912 10908
rect 8848 10848 8912 10852
rect 8928 10908 8992 10912
rect 8928 10852 8932 10908
rect 8932 10852 8988 10908
rect 8988 10852 8992 10908
rect 8928 10848 8992 10852
rect 9008 10908 9072 10912
rect 9008 10852 9012 10908
rect 9012 10852 9068 10908
rect 9068 10852 9072 10908
rect 9008 10848 9072 10852
rect 9088 10908 9152 10912
rect 9088 10852 9092 10908
rect 9092 10852 9148 10908
rect 9148 10852 9152 10908
rect 9088 10848 9152 10852
rect 11836 10780 11900 10844
rect 14412 11052 14476 11116
rect 15884 11052 15948 11116
rect 12796 10908 12860 10912
rect 12796 10852 12800 10908
rect 12800 10852 12856 10908
rect 12856 10852 12860 10908
rect 12796 10848 12860 10852
rect 12876 10908 12940 10912
rect 12876 10852 12880 10908
rect 12880 10852 12936 10908
rect 12936 10852 12940 10908
rect 12876 10848 12940 10852
rect 12956 10908 13020 10912
rect 12956 10852 12960 10908
rect 12960 10852 13016 10908
rect 13016 10852 13020 10908
rect 12956 10848 13020 10852
rect 13036 10908 13100 10912
rect 13036 10852 13040 10908
rect 13040 10852 13096 10908
rect 13096 10852 13100 10908
rect 13036 10848 13100 10852
rect 14044 10780 14108 10844
rect 15700 10780 15764 10844
rect 1900 10644 1964 10708
rect 9444 10644 9508 10708
rect 9996 10644 10060 10708
rect 10364 10644 10428 10708
rect 5580 10508 5644 10572
rect 6132 10508 6196 10572
rect 2926 10364 2990 10368
rect 2926 10308 2930 10364
rect 2930 10308 2986 10364
rect 2986 10308 2990 10364
rect 2926 10304 2990 10308
rect 3006 10364 3070 10368
rect 3006 10308 3010 10364
rect 3010 10308 3066 10364
rect 3066 10308 3070 10364
rect 3006 10304 3070 10308
rect 3086 10364 3150 10368
rect 3086 10308 3090 10364
rect 3090 10308 3146 10364
rect 3146 10308 3150 10364
rect 3086 10304 3150 10308
rect 3166 10364 3230 10368
rect 3166 10308 3170 10364
rect 3170 10308 3226 10364
rect 3226 10308 3230 10364
rect 3166 10304 3230 10308
rect 4108 10372 4172 10436
rect 7788 10508 7852 10572
rect 9444 10372 9508 10436
rect 10180 10372 10244 10436
rect 11468 10372 11532 10436
rect 12020 10508 12084 10572
rect 14596 10372 14660 10436
rect 6874 10364 6938 10368
rect 6874 10308 6878 10364
rect 6878 10308 6934 10364
rect 6934 10308 6938 10364
rect 6874 10304 6938 10308
rect 6954 10364 7018 10368
rect 6954 10308 6958 10364
rect 6958 10308 7014 10364
rect 7014 10308 7018 10364
rect 6954 10304 7018 10308
rect 7034 10364 7098 10368
rect 7034 10308 7038 10364
rect 7038 10308 7094 10364
rect 7094 10308 7098 10364
rect 7034 10304 7098 10308
rect 7114 10364 7178 10368
rect 7114 10308 7118 10364
rect 7118 10308 7174 10364
rect 7174 10308 7178 10364
rect 7114 10304 7178 10308
rect 10822 10364 10886 10368
rect 10822 10308 10826 10364
rect 10826 10308 10882 10364
rect 10882 10308 10886 10364
rect 10822 10304 10886 10308
rect 10902 10364 10966 10368
rect 10902 10308 10906 10364
rect 10906 10308 10962 10364
rect 10962 10308 10966 10364
rect 10902 10304 10966 10308
rect 10982 10364 11046 10368
rect 10982 10308 10986 10364
rect 10986 10308 11042 10364
rect 11042 10308 11046 10364
rect 10982 10304 11046 10308
rect 11062 10364 11126 10368
rect 11062 10308 11066 10364
rect 11066 10308 11122 10364
rect 11122 10308 11126 10364
rect 11062 10304 11126 10308
rect 14770 10364 14834 10368
rect 14770 10308 14774 10364
rect 14774 10308 14830 10364
rect 14830 10308 14834 10364
rect 14770 10304 14834 10308
rect 14850 10364 14914 10368
rect 14850 10308 14854 10364
rect 14854 10308 14910 10364
rect 14910 10308 14914 10364
rect 14850 10304 14914 10308
rect 14930 10364 14994 10368
rect 14930 10308 14934 10364
rect 14934 10308 14990 10364
rect 14990 10308 14994 10364
rect 14930 10304 14994 10308
rect 15010 10364 15074 10368
rect 15010 10308 15014 10364
rect 15014 10308 15070 10364
rect 15070 10308 15074 10364
rect 15010 10304 15074 10308
rect 4292 10100 4356 10164
rect 6132 9828 6196 9892
rect 8524 10100 8588 10164
rect 9996 9964 10060 10028
rect 16436 9828 16500 9892
rect 4900 9820 4964 9824
rect 4900 9764 4904 9820
rect 4904 9764 4960 9820
rect 4960 9764 4964 9820
rect 4900 9760 4964 9764
rect 4980 9820 5044 9824
rect 4980 9764 4984 9820
rect 4984 9764 5040 9820
rect 5040 9764 5044 9820
rect 4980 9760 5044 9764
rect 5060 9820 5124 9824
rect 5060 9764 5064 9820
rect 5064 9764 5120 9820
rect 5120 9764 5124 9820
rect 5060 9760 5124 9764
rect 5140 9820 5204 9824
rect 5140 9764 5144 9820
rect 5144 9764 5200 9820
rect 5200 9764 5204 9820
rect 5140 9760 5204 9764
rect 8848 9820 8912 9824
rect 8848 9764 8852 9820
rect 8852 9764 8908 9820
rect 8908 9764 8912 9820
rect 8848 9760 8912 9764
rect 8928 9820 8992 9824
rect 8928 9764 8932 9820
rect 8932 9764 8988 9820
rect 8988 9764 8992 9820
rect 8928 9760 8992 9764
rect 9008 9820 9072 9824
rect 9008 9764 9012 9820
rect 9012 9764 9068 9820
rect 9068 9764 9072 9820
rect 9008 9760 9072 9764
rect 9088 9820 9152 9824
rect 9088 9764 9092 9820
rect 9092 9764 9148 9820
rect 9148 9764 9152 9820
rect 9088 9760 9152 9764
rect 12796 9820 12860 9824
rect 12796 9764 12800 9820
rect 12800 9764 12856 9820
rect 12856 9764 12860 9820
rect 12796 9760 12860 9764
rect 12876 9820 12940 9824
rect 12876 9764 12880 9820
rect 12880 9764 12936 9820
rect 12936 9764 12940 9820
rect 12876 9760 12940 9764
rect 12956 9820 13020 9824
rect 12956 9764 12960 9820
rect 12960 9764 13016 9820
rect 13016 9764 13020 9820
rect 12956 9760 13020 9764
rect 13036 9820 13100 9824
rect 13036 9764 13040 9820
rect 13040 9764 13096 9820
rect 13096 9764 13100 9820
rect 13036 9760 13100 9764
rect 7604 9692 7668 9756
rect 9628 9752 9692 9756
rect 9628 9696 9642 9752
rect 9642 9696 9692 9752
rect 9628 9692 9692 9696
rect 10180 9692 10244 9756
rect 11284 9556 11348 9620
rect 11652 9556 11716 9620
rect 3740 9420 3804 9484
rect 10548 9420 10612 9484
rect 13308 9420 13372 9484
rect 6684 9284 6748 9348
rect 2926 9276 2990 9280
rect 2926 9220 2930 9276
rect 2930 9220 2986 9276
rect 2986 9220 2990 9276
rect 2926 9216 2990 9220
rect 3006 9276 3070 9280
rect 3006 9220 3010 9276
rect 3010 9220 3066 9276
rect 3066 9220 3070 9276
rect 3006 9216 3070 9220
rect 3086 9276 3150 9280
rect 3086 9220 3090 9276
rect 3090 9220 3146 9276
rect 3146 9220 3150 9276
rect 3086 9216 3150 9220
rect 3166 9276 3230 9280
rect 3166 9220 3170 9276
rect 3170 9220 3226 9276
rect 3226 9220 3230 9276
rect 3166 9216 3230 9220
rect 6874 9276 6938 9280
rect 6874 9220 6878 9276
rect 6878 9220 6934 9276
rect 6934 9220 6938 9276
rect 6874 9216 6938 9220
rect 6954 9276 7018 9280
rect 6954 9220 6958 9276
rect 6958 9220 7014 9276
rect 7014 9220 7018 9276
rect 6954 9216 7018 9220
rect 7034 9276 7098 9280
rect 7034 9220 7038 9276
rect 7038 9220 7094 9276
rect 7094 9220 7098 9276
rect 7034 9216 7098 9220
rect 7114 9276 7178 9280
rect 7114 9220 7118 9276
rect 7118 9220 7174 9276
rect 7174 9220 7178 9276
rect 7114 9216 7178 9220
rect 10822 9276 10886 9280
rect 10822 9220 10826 9276
rect 10826 9220 10882 9276
rect 10882 9220 10886 9276
rect 10822 9216 10886 9220
rect 10902 9276 10966 9280
rect 10902 9220 10906 9276
rect 10906 9220 10962 9276
rect 10962 9220 10966 9276
rect 10902 9216 10966 9220
rect 10982 9276 11046 9280
rect 10982 9220 10986 9276
rect 10986 9220 11042 9276
rect 11042 9220 11046 9276
rect 10982 9216 11046 9220
rect 11062 9276 11126 9280
rect 11062 9220 11066 9276
rect 11066 9220 11122 9276
rect 11122 9220 11126 9276
rect 11062 9216 11126 9220
rect 14770 9276 14834 9280
rect 14770 9220 14774 9276
rect 14774 9220 14830 9276
rect 14830 9220 14834 9276
rect 14770 9216 14834 9220
rect 14850 9276 14914 9280
rect 14850 9220 14854 9276
rect 14854 9220 14910 9276
rect 14910 9220 14914 9276
rect 14850 9216 14914 9220
rect 14930 9276 14994 9280
rect 14930 9220 14934 9276
rect 14934 9220 14990 9276
rect 14990 9220 14994 9276
rect 14930 9216 14994 9220
rect 15010 9276 15074 9280
rect 15010 9220 15014 9276
rect 15014 9220 15070 9276
rect 15070 9220 15074 9276
rect 15010 9216 15074 9220
rect 14044 9072 14108 9076
rect 14044 9016 14058 9072
rect 14058 9016 14108 9072
rect 14044 9012 14108 9016
rect 15700 9012 15764 9076
rect 10548 8740 10612 8804
rect 13860 8876 13924 8940
rect 4900 8732 4964 8736
rect 4900 8676 4904 8732
rect 4904 8676 4960 8732
rect 4960 8676 4964 8732
rect 4900 8672 4964 8676
rect 4980 8732 5044 8736
rect 4980 8676 4984 8732
rect 4984 8676 5040 8732
rect 5040 8676 5044 8732
rect 4980 8672 5044 8676
rect 5060 8732 5124 8736
rect 5060 8676 5064 8732
rect 5064 8676 5120 8732
rect 5120 8676 5124 8732
rect 5060 8672 5124 8676
rect 5140 8732 5204 8736
rect 5140 8676 5144 8732
rect 5144 8676 5200 8732
rect 5200 8676 5204 8732
rect 5140 8672 5204 8676
rect 8848 8732 8912 8736
rect 8848 8676 8852 8732
rect 8852 8676 8908 8732
rect 8908 8676 8912 8732
rect 8848 8672 8912 8676
rect 8928 8732 8992 8736
rect 8928 8676 8932 8732
rect 8932 8676 8988 8732
rect 8988 8676 8992 8732
rect 8928 8672 8992 8676
rect 9008 8732 9072 8736
rect 9008 8676 9012 8732
rect 9012 8676 9068 8732
rect 9068 8676 9072 8732
rect 9008 8672 9072 8676
rect 9088 8732 9152 8736
rect 9088 8676 9092 8732
rect 9092 8676 9148 8732
rect 9148 8676 9152 8732
rect 9088 8672 9152 8676
rect 12796 8732 12860 8736
rect 12796 8676 12800 8732
rect 12800 8676 12856 8732
rect 12856 8676 12860 8732
rect 12796 8672 12860 8676
rect 12876 8732 12940 8736
rect 12876 8676 12880 8732
rect 12880 8676 12936 8732
rect 12936 8676 12940 8732
rect 12876 8672 12940 8676
rect 12956 8732 13020 8736
rect 12956 8676 12960 8732
rect 12960 8676 13016 8732
rect 13016 8676 13020 8732
rect 12956 8672 13020 8676
rect 13036 8732 13100 8736
rect 13036 8676 13040 8732
rect 13040 8676 13096 8732
rect 13096 8676 13100 8732
rect 13036 8672 13100 8676
rect 12572 8664 12636 8668
rect 12572 8608 12586 8664
rect 12586 8608 12636 8664
rect 12572 8604 12636 8608
rect 13308 8604 13372 8668
rect 14412 8604 14476 8668
rect 4476 8332 4540 8396
rect 4660 8332 4724 8396
rect 14412 8468 14476 8532
rect 11652 8332 11716 8396
rect 12204 8332 12268 8396
rect 16068 8468 16132 8532
rect 15700 8392 15764 8396
rect 15700 8336 15750 8392
rect 15750 8336 15764 8392
rect 15700 8332 15764 8336
rect 8156 8196 8220 8260
rect 9628 8196 9692 8260
rect 14228 8196 14292 8260
rect 2926 8188 2990 8192
rect 2926 8132 2930 8188
rect 2930 8132 2986 8188
rect 2986 8132 2990 8188
rect 2926 8128 2990 8132
rect 3006 8188 3070 8192
rect 3006 8132 3010 8188
rect 3010 8132 3066 8188
rect 3066 8132 3070 8188
rect 3006 8128 3070 8132
rect 3086 8188 3150 8192
rect 3086 8132 3090 8188
rect 3090 8132 3146 8188
rect 3146 8132 3150 8188
rect 3086 8128 3150 8132
rect 3166 8188 3230 8192
rect 3166 8132 3170 8188
rect 3170 8132 3226 8188
rect 3226 8132 3230 8188
rect 3166 8128 3230 8132
rect 6874 8188 6938 8192
rect 6874 8132 6878 8188
rect 6878 8132 6934 8188
rect 6934 8132 6938 8188
rect 6874 8128 6938 8132
rect 6954 8188 7018 8192
rect 6954 8132 6958 8188
rect 6958 8132 7014 8188
rect 7014 8132 7018 8188
rect 6954 8128 7018 8132
rect 7034 8188 7098 8192
rect 7034 8132 7038 8188
rect 7038 8132 7094 8188
rect 7094 8132 7098 8188
rect 7034 8128 7098 8132
rect 7114 8188 7178 8192
rect 7114 8132 7118 8188
rect 7118 8132 7174 8188
rect 7174 8132 7178 8188
rect 7114 8128 7178 8132
rect 10822 8188 10886 8192
rect 10822 8132 10826 8188
rect 10826 8132 10882 8188
rect 10882 8132 10886 8188
rect 10822 8128 10886 8132
rect 10902 8188 10966 8192
rect 10902 8132 10906 8188
rect 10906 8132 10962 8188
rect 10962 8132 10966 8188
rect 10902 8128 10966 8132
rect 10982 8188 11046 8192
rect 10982 8132 10986 8188
rect 10986 8132 11042 8188
rect 11042 8132 11046 8188
rect 10982 8128 11046 8132
rect 11062 8188 11126 8192
rect 11062 8132 11066 8188
rect 11066 8132 11122 8188
rect 11122 8132 11126 8188
rect 11062 8128 11126 8132
rect 14770 8188 14834 8192
rect 14770 8132 14774 8188
rect 14774 8132 14830 8188
rect 14830 8132 14834 8188
rect 14770 8128 14834 8132
rect 14850 8188 14914 8192
rect 14850 8132 14854 8188
rect 14854 8132 14910 8188
rect 14910 8132 14914 8188
rect 14850 8128 14914 8132
rect 14930 8188 14994 8192
rect 14930 8132 14934 8188
rect 14934 8132 14990 8188
rect 14990 8132 14994 8188
rect 14930 8128 14994 8132
rect 15010 8188 15074 8192
rect 15010 8132 15014 8188
rect 15014 8132 15070 8188
rect 15070 8132 15074 8188
rect 15010 8128 15074 8132
rect 7604 8060 7668 8124
rect 9812 8060 9876 8124
rect 5764 7924 5828 7988
rect 9628 7924 9692 7988
rect 11836 8060 11900 8124
rect 12388 8060 12452 8124
rect 4292 7788 4356 7852
rect 5580 7652 5644 7716
rect 4900 7644 4964 7648
rect 4900 7588 4904 7644
rect 4904 7588 4960 7644
rect 4960 7588 4964 7644
rect 4900 7584 4964 7588
rect 4980 7644 5044 7648
rect 4980 7588 4984 7644
rect 4984 7588 5040 7644
rect 5040 7588 5044 7644
rect 4980 7584 5044 7588
rect 5060 7644 5124 7648
rect 5060 7588 5064 7644
rect 5064 7588 5120 7644
rect 5120 7588 5124 7644
rect 5060 7584 5124 7588
rect 5140 7644 5204 7648
rect 5140 7588 5144 7644
rect 5144 7588 5200 7644
rect 5200 7588 5204 7644
rect 5140 7584 5204 7588
rect 8848 7644 8912 7648
rect 8848 7588 8852 7644
rect 8852 7588 8908 7644
rect 8908 7588 8912 7644
rect 8848 7584 8912 7588
rect 8928 7644 8992 7648
rect 8928 7588 8932 7644
rect 8932 7588 8988 7644
rect 8988 7588 8992 7644
rect 8928 7584 8992 7588
rect 9008 7644 9072 7648
rect 9008 7588 9012 7644
rect 9012 7588 9068 7644
rect 9068 7588 9072 7644
rect 9008 7584 9072 7588
rect 9088 7644 9152 7648
rect 9088 7588 9092 7644
rect 9092 7588 9148 7644
rect 9148 7588 9152 7644
rect 9088 7584 9152 7588
rect 9628 7788 9692 7852
rect 12388 7924 12452 7988
rect 11468 7848 11532 7852
rect 11468 7792 11482 7848
rect 11482 7792 11532 7848
rect 11468 7788 11532 7792
rect 12204 7788 12268 7852
rect 12572 7788 12636 7852
rect 13860 7848 13924 7852
rect 13860 7792 13874 7848
rect 13874 7792 13924 7848
rect 13860 7788 13924 7792
rect 9444 7652 9508 7716
rect 12796 7644 12860 7648
rect 12796 7588 12800 7644
rect 12800 7588 12856 7644
rect 12856 7588 12860 7644
rect 12796 7584 12860 7588
rect 12876 7644 12940 7648
rect 12876 7588 12880 7644
rect 12880 7588 12936 7644
rect 12936 7588 12940 7644
rect 12876 7584 12940 7588
rect 12956 7644 13020 7648
rect 12956 7588 12960 7644
rect 12960 7588 13016 7644
rect 13016 7588 13020 7644
rect 12956 7584 13020 7588
rect 13036 7644 13100 7648
rect 13036 7588 13040 7644
rect 13040 7588 13096 7644
rect 13096 7588 13100 7644
rect 13036 7584 13100 7588
rect 4108 7380 4172 7444
rect 9996 7380 10060 7444
rect 16620 7516 16684 7580
rect 9812 7168 9876 7172
rect 9812 7112 9826 7168
rect 9826 7112 9876 7168
rect 9812 7108 9876 7112
rect 11284 7108 11348 7172
rect 2926 7100 2990 7104
rect 2926 7044 2930 7100
rect 2930 7044 2986 7100
rect 2986 7044 2990 7100
rect 2926 7040 2990 7044
rect 3006 7100 3070 7104
rect 3006 7044 3010 7100
rect 3010 7044 3066 7100
rect 3066 7044 3070 7100
rect 3006 7040 3070 7044
rect 3086 7100 3150 7104
rect 3086 7044 3090 7100
rect 3090 7044 3146 7100
rect 3146 7044 3150 7100
rect 3086 7040 3150 7044
rect 3166 7100 3230 7104
rect 3166 7044 3170 7100
rect 3170 7044 3226 7100
rect 3226 7044 3230 7100
rect 3166 7040 3230 7044
rect 6874 7100 6938 7104
rect 6874 7044 6878 7100
rect 6878 7044 6934 7100
rect 6934 7044 6938 7100
rect 6874 7040 6938 7044
rect 6954 7100 7018 7104
rect 6954 7044 6958 7100
rect 6958 7044 7014 7100
rect 7014 7044 7018 7100
rect 6954 7040 7018 7044
rect 7034 7100 7098 7104
rect 7034 7044 7038 7100
rect 7038 7044 7094 7100
rect 7094 7044 7098 7100
rect 7034 7040 7098 7044
rect 7114 7100 7178 7104
rect 7114 7044 7118 7100
rect 7118 7044 7174 7100
rect 7174 7044 7178 7100
rect 7114 7040 7178 7044
rect 10822 7100 10886 7104
rect 10822 7044 10826 7100
rect 10826 7044 10882 7100
rect 10882 7044 10886 7100
rect 10822 7040 10886 7044
rect 10902 7100 10966 7104
rect 10902 7044 10906 7100
rect 10906 7044 10962 7100
rect 10962 7044 10966 7100
rect 10902 7040 10966 7044
rect 10982 7100 11046 7104
rect 10982 7044 10986 7100
rect 10986 7044 11042 7100
rect 11042 7044 11046 7100
rect 10982 7040 11046 7044
rect 11062 7100 11126 7104
rect 11062 7044 11066 7100
rect 11066 7044 11122 7100
rect 11122 7044 11126 7100
rect 11062 7040 11126 7044
rect 14770 7100 14834 7104
rect 14770 7044 14774 7100
rect 14774 7044 14830 7100
rect 14830 7044 14834 7100
rect 14770 7040 14834 7044
rect 14850 7100 14914 7104
rect 14850 7044 14854 7100
rect 14854 7044 14910 7100
rect 14910 7044 14914 7100
rect 14850 7040 14914 7044
rect 14930 7100 14994 7104
rect 14930 7044 14934 7100
rect 14934 7044 14990 7100
rect 14990 7044 14994 7100
rect 14930 7040 14994 7044
rect 15010 7100 15074 7104
rect 15010 7044 15014 7100
rect 15014 7044 15070 7100
rect 15070 7044 15074 7100
rect 15010 7040 15074 7044
rect 9260 6972 9324 7036
rect 2636 6896 2700 6900
rect 2636 6840 2686 6896
rect 2686 6840 2700 6896
rect 2636 6836 2700 6840
rect 11284 6836 11348 6900
rect 15332 6836 15396 6900
rect 10180 6700 10244 6764
rect 15332 6564 15396 6628
rect 15700 6564 15764 6628
rect 4900 6556 4964 6560
rect 4900 6500 4904 6556
rect 4904 6500 4960 6556
rect 4960 6500 4964 6556
rect 4900 6496 4964 6500
rect 4980 6556 5044 6560
rect 4980 6500 4984 6556
rect 4984 6500 5040 6556
rect 5040 6500 5044 6556
rect 4980 6496 5044 6500
rect 5060 6556 5124 6560
rect 5060 6500 5064 6556
rect 5064 6500 5120 6556
rect 5120 6500 5124 6556
rect 5060 6496 5124 6500
rect 5140 6556 5204 6560
rect 5140 6500 5144 6556
rect 5144 6500 5200 6556
rect 5200 6500 5204 6556
rect 5140 6496 5204 6500
rect 8848 6556 8912 6560
rect 8848 6500 8852 6556
rect 8852 6500 8908 6556
rect 8908 6500 8912 6556
rect 8848 6496 8912 6500
rect 8928 6556 8992 6560
rect 8928 6500 8932 6556
rect 8932 6500 8988 6556
rect 8988 6500 8992 6556
rect 8928 6496 8992 6500
rect 9008 6556 9072 6560
rect 9008 6500 9012 6556
rect 9012 6500 9068 6556
rect 9068 6500 9072 6556
rect 9008 6496 9072 6500
rect 9088 6556 9152 6560
rect 9088 6500 9092 6556
rect 9092 6500 9148 6556
rect 9148 6500 9152 6556
rect 9088 6496 9152 6500
rect 12796 6556 12860 6560
rect 12796 6500 12800 6556
rect 12800 6500 12856 6556
rect 12856 6500 12860 6556
rect 12796 6496 12860 6500
rect 12876 6556 12940 6560
rect 12876 6500 12880 6556
rect 12880 6500 12936 6556
rect 12936 6500 12940 6556
rect 12876 6496 12940 6500
rect 12956 6556 13020 6560
rect 12956 6500 12960 6556
rect 12960 6500 13016 6556
rect 13016 6500 13020 6556
rect 12956 6496 13020 6500
rect 13036 6556 13100 6560
rect 13036 6500 13040 6556
rect 13040 6500 13096 6556
rect 13096 6500 13100 6556
rect 13036 6496 13100 6500
rect 8156 6488 8220 6492
rect 8156 6432 8206 6488
rect 8206 6432 8220 6488
rect 8156 6428 8220 6432
rect 13676 6428 13740 6492
rect 8524 6292 8588 6356
rect 12388 6292 12452 6356
rect 13860 6292 13924 6356
rect 16252 6156 16316 6220
rect 2926 6012 2990 6016
rect 2926 5956 2930 6012
rect 2930 5956 2986 6012
rect 2986 5956 2990 6012
rect 2926 5952 2990 5956
rect 3006 6012 3070 6016
rect 3006 5956 3010 6012
rect 3010 5956 3066 6012
rect 3066 5956 3070 6012
rect 3006 5952 3070 5956
rect 3086 6012 3150 6016
rect 3086 5956 3090 6012
rect 3090 5956 3146 6012
rect 3146 5956 3150 6012
rect 3086 5952 3150 5956
rect 3166 6012 3230 6016
rect 3166 5956 3170 6012
rect 3170 5956 3226 6012
rect 3226 5956 3230 6012
rect 3166 5952 3230 5956
rect 6874 6012 6938 6016
rect 6874 5956 6878 6012
rect 6878 5956 6934 6012
rect 6934 5956 6938 6012
rect 6874 5952 6938 5956
rect 6954 6012 7018 6016
rect 6954 5956 6958 6012
rect 6958 5956 7014 6012
rect 7014 5956 7018 6012
rect 6954 5952 7018 5956
rect 7034 6012 7098 6016
rect 7034 5956 7038 6012
rect 7038 5956 7094 6012
rect 7094 5956 7098 6012
rect 7034 5952 7098 5956
rect 7114 6012 7178 6016
rect 7114 5956 7118 6012
rect 7118 5956 7174 6012
rect 7174 5956 7178 6012
rect 7114 5952 7178 5956
rect 4108 5672 4172 5676
rect 4108 5616 4122 5672
rect 4122 5616 4172 5672
rect 4108 5612 4172 5616
rect 6316 5748 6380 5812
rect 9628 5884 9692 5948
rect 11468 6020 11532 6084
rect 10822 6012 10886 6016
rect 10822 5956 10826 6012
rect 10826 5956 10882 6012
rect 10882 5956 10886 6012
rect 10822 5952 10886 5956
rect 10902 6012 10966 6016
rect 10902 5956 10906 6012
rect 10906 5956 10962 6012
rect 10962 5956 10966 6012
rect 10902 5952 10966 5956
rect 10982 6012 11046 6016
rect 10982 5956 10986 6012
rect 10986 5956 11042 6012
rect 11042 5956 11046 6012
rect 10982 5952 11046 5956
rect 11062 6012 11126 6016
rect 11062 5956 11066 6012
rect 11066 5956 11122 6012
rect 11122 5956 11126 6012
rect 11062 5952 11126 5956
rect 14770 6012 14834 6016
rect 14770 5956 14774 6012
rect 14774 5956 14830 6012
rect 14830 5956 14834 6012
rect 14770 5952 14834 5956
rect 14850 6012 14914 6016
rect 14850 5956 14854 6012
rect 14854 5956 14910 6012
rect 14910 5956 14914 6012
rect 14850 5952 14914 5956
rect 14930 6012 14994 6016
rect 14930 5956 14934 6012
rect 14934 5956 14990 6012
rect 14990 5956 14994 6012
rect 14930 5952 14994 5956
rect 15010 6012 15074 6016
rect 15010 5956 15014 6012
rect 15014 5956 15070 6012
rect 15070 5956 15074 6012
rect 15010 5952 15074 5956
rect 14412 5884 14476 5948
rect 13676 5748 13740 5812
rect 9628 5476 9692 5540
rect 10364 5476 10428 5540
rect 11468 5476 11532 5540
rect 4900 5468 4964 5472
rect 4900 5412 4904 5468
rect 4904 5412 4960 5468
rect 4960 5412 4964 5468
rect 4900 5408 4964 5412
rect 4980 5468 5044 5472
rect 4980 5412 4984 5468
rect 4984 5412 5040 5468
rect 5040 5412 5044 5468
rect 4980 5408 5044 5412
rect 5060 5468 5124 5472
rect 5060 5412 5064 5468
rect 5064 5412 5120 5468
rect 5120 5412 5124 5468
rect 5060 5408 5124 5412
rect 5140 5468 5204 5472
rect 5140 5412 5144 5468
rect 5144 5412 5200 5468
rect 5200 5412 5204 5468
rect 5140 5408 5204 5412
rect 8848 5468 8912 5472
rect 8848 5412 8852 5468
rect 8852 5412 8908 5468
rect 8908 5412 8912 5468
rect 8848 5408 8912 5412
rect 8928 5468 8992 5472
rect 8928 5412 8932 5468
rect 8932 5412 8988 5468
rect 8988 5412 8992 5468
rect 8928 5408 8992 5412
rect 9008 5468 9072 5472
rect 9008 5412 9012 5468
rect 9012 5412 9068 5468
rect 9068 5412 9072 5468
rect 9008 5408 9072 5412
rect 9088 5468 9152 5472
rect 9088 5412 9092 5468
rect 9092 5412 9148 5468
rect 9148 5412 9152 5468
rect 9088 5408 9152 5412
rect 7972 5340 8036 5404
rect 9260 5340 9324 5404
rect 12204 5476 12268 5540
rect 12796 5468 12860 5472
rect 12796 5412 12800 5468
rect 12800 5412 12856 5468
rect 12856 5412 12860 5468
rect 12796 5408 12860 5412
rect 12876 5468 12940 5472
rect 12876 5412 12880 5468
rect 12880 5412 12936 5468
rect 12936 5412 12940 5468
rect 12876 5408 12940 5412
rect 12956 5468 13020 5472
rect 12956 5412 12960 5468
rect 12960 5412 13016 5468
rect 13016 5412 13020 5468
rect 12956 5408 13020 5412
rect 13036 5468 13100 5472
rect 13036 5412 13040 5468
rect 13040 5412 13096 5468
rect 13096 5412 13100 5468
rect 13036 5408 13100 5412
rect 6684 5204 6748 5268
rect 6132 5068 6196 5132
rect 15148 5068 15212 5132
rect 10364 4932 10428 4996
rect 12020 4932 12084 4996
rect 12204 4932 12268 4996
rect 2926 4924 2990 4928
rect 2926 4868 2930 4924
rect 2930 4868 2986 4924
rect 2986 4868 2990 4924
rect 2926 4864 2990 4868
rect 3006 4924 3070 4928
rect 3006 4868 3010 4924
rect 3010 4868 3066 4924
rect 3066 4868 3070 4924
rect 3006 4864 3070 4868
rect 3086 4924 3150 4928
rect 3086 4868 3090 4924
rect 3090 4868 3146 4924
rect 3146 4868 3150 4924
rect 3086 4864 3150 4868
rect 3166 4924 3230 4928
rect 3166 4868 3170 4924
rect 3170 4868 3226 4924
rect 3226 4868 3230 4924
rect 3166 4864 3230 4868
rect 6874 4924 6938 4928
rect 6874 4868 6878 4924
rect 6878 4868 6934 4924
rect 6934 4868 6938 4924
rect 6874 4864 6938 4868
rect 6954 4924 7018 4928
rect 6954 4868 6958 4924
rect 6958 4868 7014 4924
rect 7014 4868 7018 4924
rect 6954 4864 7018 4868
rect 7034 4924 7098 4928
rect 7034 4868 7038 4924
rect 7038 4868 7094 4924
rect 7094 4868 7098 4924
rect 7034 4864 7098 4868
rect 7114 4924 7178 4928
rect 7114 4868 7118 4924
rect 7118 4868 7174 4924
rect 7174 4868 7178 4924
rect 7114 4864 7178 4868
rect 10822 4924 10886 4928
rect 10822 4868 10826 4924
rect 10826 4868 10882 4924
rect 10882 4868 10886 4924
rect 10822 4864 10886 4868
rect 10902 4924 10966 4928
rect 10902 4868 10906 4924
rect 10906 4868 10962 4924
rect 10962 4868 10966 4924
rect 10902 4864 10966 4868
rect 10982 4924 11046 4928
rect 10982 4868 10986 4924
rect 10986 4868 11042 4924
rect 11042 4868 11046 4924
rect 10982 4864 11046 4868
rect 11062 4924 11126 4928
rect 11062 4868 11066 4924
rect 11066 4868 11122 4924
rect 11122 4868 11126 4924
rect 11062 4864 11126 4868
rect 14770 4924 14834 4928
rect 14770 4868 14774 4924
rect 14774 4868 14830 4924
rect 14830 4868 14834 4924
rect 14770 4864 14834 4868
rect 14850 4924 14914 4928
rect 14850 4868 14854 4924
rect 14854 4868 14910 4924
rect 14910 4868 14914 4924
rect 14850 4864 14914 4868
rect 14930 4924 14994 4928
rect 14930 4868 14934 4924
rect 14934 4868 14990 4924
rect 14990 4868 14994 4924
rect 14930 4864 14994 4868
rect 15010 4924 15074 4928
rect 15010 4868 15014 4924
rect 15014 4868 15070 4924
rect 15070 4868 15074 4924
rect 15010 4864 15074 4868
rect 8708 4796 8772 4860
rect 9812 4796 9876 4860
rect 11836 4796 11900 4860
rect 9628 4720 9692 4724
rect 9628 4664 9678 4720
rect 9678 4664 9692 4720
rect 7788 4524 7852 4588
rect 9628 4660 9692 4664
rect 9812 4660 9876 4724
rect 11284 4660 11348 4724
rect 13492 4796 13556 4860
rect 12020 4660 12084 4724
rect 13308 4660 13372 4724
rect 4900 4380 4964 4384
rect 4900 4324 4904 4380
rect 4904 4324 4960 4380
rect 4960 4324 4964 4380
rect 4900 4320 4964 4324
rect 4980 4380 5044 4384
rect 4980 4324 4984 4380
rect 4984 4324 5040 4380
rect 5040 4324 5044 4380
rect 4980 4320 5044 4324
rect 5060 4380 5124 4384
rect 5060 4324 5064 4380
rect 5064 4324 5120 4380
rect 5120 4324 5124 4380
rect 5060 4320 5124 4324
rect 5140 4380 5204 4384
rect 5140 4324 5144 4380
rect 5144 4324 5200 4380
rect 5200 4324 5204 4380
rect 5140 4320 5204 4324
rect 14228 4388 14292 4452
rect 8848 4380 8912 4384
rect 8848 4324 8852 4380
rect 8852 4324 8908 4380
rect 8908 4324 8912 4380
rect 8848 4320 8912 4324
rect 8928 4380 8992 4384
rect 8928 4324 8932 4380
rect 8932 4324 8988 4380
rect 8988 4324 8992 4380
rect 8928 4320 8992 4324
rect 9008 4380 9072 4384
rect 9008 4324 9012 4380
rect 9012 4324 9068 4380
rect 9068 4324 9072 4380
rect 9008 4320 9072 4324
rect 9088 4380 9152 4384
rect 9088 4324 9092 4380
rect 9092 4324 9148 4380
rect 9148 4324 9152 4380
rect 9088 4320 9152 4324
rect 12796 4380 12860 4384
rect 12796 4324 12800 4380
rect 12800 4324 12856 4380
rect 12856 4324 12860 4380
rect 12796 4320 12860 4324
rect 12876 4380 12940 4384
rect 12876 4324 12880 4380
rect 12880 4324 12936 4380
rect 12936 4324 12940 4380
rect 12876 4320 12940 4324
rect 12956 4380 13020 4384
rect 12956 4324 12960 4380
rect 12960 4324 13016 4380
rect 13016 4324 13020 4380
rect 12956 4320 13020 4324
rect 13036 4380 13100 4384
rect 13036 4324 13040 4380
rect 13040 4324 13096 4380
rect 13096 4324 13100 4380
rect 13036 4320 13100 4324
rect 8708 4252 8772 4316
rect 7972 4116 8036 4180
rect 15516 4116 15580 4180
rect 16804 4116 16868 4180
rect 6316 3844 6380 3908
rect 7420 3904 7484 3908
rect 7420 3848 7434 3904
rect 7434 3848 7484 3904
rect 7420 3844 7484 3848
rect 7788 3844 7852 3908
rect 9996 3844 10060 3908
rect 12020 3844 12084 3908
rect 2926 3836 2990 3840
rect 2926 3780 2930 3836
rect 2930 3780 2986 3836
rect 2986 3780 2990 3836
rect 2926 3776 2990 3780
rect 3006 3836 3070 3840
rect 3006 3780 3010 3836
rect 3010 3780 3066 3836
rect 3066 3780 3070 3836
rect 3006 3776 3070 3780
rect 3086 3836 3150 3840
rect 3086 3780 3090 3836
rect 3090 3780 3146 3836
rect 3146 3780 3150 3836
rect 3086 3776 3150 3780
rect 3166 3836 3230 3840
rect 3166 3780 3170 3836
rect 3170 3780 3226 3836
rect 3226 3780 3230 3836
rect 3166 3776 3230 3780
rect 6874 3836 6938 3840
rect 6874 3780 6878 3836
rect 6878 3780 6934 3836
rect 6934 3780 6938 3836
rect 6874 3776 6938 3780
rect 6954 3836 7018 3840
rect 6954 3780 6958 3836
rect 6958 3780 7014 3836
rect 7014 3780 7018 3836
rect 6954 3776 7018 3780
rect 7034 3836 7098 3840
rect 7034 3780 7038 3836
rect 7038 3780 7094 3836
rect 7094 3780 7098 3836
rect 7034 3776 7098 3780
rect 7114 3836 7178 3840
rect 7114 3780 7118 3836
rect 7118 3780 7174 3836
rect 7174 3780 7178 3836
rect 7114 3776 7178 3780
rect 10822 3836 10886 3840
rect 10822 3780 10826 3836
rect 10826 3780 10882 3836
rect 10882 3780 10886 3836
rect 10822 3776 10886 3780
rect 10902 3836 10966 3840
rect 10902 3780 10906 3836
rect 10906 3780 10962 3836
rect 10962 3780 10966 3836
rect 10902 3776 10966 3780
rect 10982 3836 11046 3840
rect 10982 3780 10986 3836
rect 10986 3780 11042 3836
rect 11042 3780 11046 3836
rect 10982 3776 11046 3780
rect 11062 3836 11126 3840
rect 11062 3780 11066 3836
rect 11066 3780 11122 3836
rect 11122 3780 11126 3836
rect 11062 3776 11126 3780
rect 14770 3836 14834 3840
rect 14770 3780 14774 3836
rect 14774 3780 14830 3836
rect 14830 3780 14834 3836
rect 14770 3776 14834 3780
rect 14850 3836 14914 3840
rect 14850 3780 14854 3836
rect 14854 3780 14910 3836
rect 14910 3780 14914 3836
rect 14850 3776 14914 3780
rect 14930 3836 14994 3840
rect 14930 3780 14934 3836
rect 14934 3780 14990 3836
rect 14990 3780 14994 3836
rect 14930 3776 14994 3780
rect 15010 3836 15074 3840
rect 15010 3780 15014 3836
rect 15014 3780 15070 3836
rect 15070 3780 15074 3836
rect 15010 3776 15074 3780
rect 5764 3768 5828 3772
rect 5764 3712 5814 3768
rect 5814 3712 5828 3768
rect 5764 3708 5828 3712
rect 8340 3708 8404 3772
rect 8708 3708 8772 3772
rect 11652 3708 11716 3772
rect 2636 3436 2700 3500
rect 7972 3496 8036 3500
rect 7972 3440 8022 3496
rect 8022 3440 8036 3496
rect 7972 3436 8036 3440
rect 14044 3572 14108 3636
rect 4292 3300 4356 3364
rect 7604 3300 7668 3364
rect 8524 3300 8588 3364
rect 4900 3292 4964 3296
rect 4900 3236 4904 3292
rect 4904 3236 4960 3292
rect 4960 3236 4964 3292
rect 4900 3232 4964 3236
rect 4980 3292 5044 3296
rect 4980 3236 4984 3292
rect 4984 3236 5040 3292
rect 5040 3236 5044 3292
rect 4980 3232 5044 3236
rect 5060 3292 5124 3296
rect 5060 3236 5064 3292
rect 5064 3236 5120 3292
rect 5120 3236 5124 3292
rect 5060 3232 5124 3236
rect 5140 3292 5204 3296
rect 5140 3236 5144 3292
rect 5144 3236 5200 3292
rect 5200 3236 5204 3292
rect 5140 3232 5204 3236
rect 5580 3164 5644 3228
rect 8848 3292 8912 3296
rect 8848 3236 8852 3292
rect 8852 3236 8908 3292
rect 8908 3236 8912 3292
rect 8848 3232 8912 3236
rect 8928 3292 8992 3296
rect 8928 3236 8932 3292
rect 8932 3236 8988 3292
rect 8988 3236 8992 3292
rect 8928 3232 8992 3236
rect 9008 3292 9072 3296
rect 9008 3236 9012 3292
rect 9012 3236 9068 3292
rect 9068 3236 9072 3292
rect 9008 3232 9072 3236
rect 9088 3292 9152 3296
rect 9088 3236 9092 3292
rect 9092 3236 9148 3292
rect 9148 3236 9152 3292
rect 9088 3232 9152 3236
rect 12796 3292 12860 3296
rect 12796 3236 12800 3292
rect 12800 3236 12856 3292
rect 12856 3236 12860 3292
rect 12796 3232 12860 3236
rect 12876 3292 12940 3296
rect 12876 3236 12880 3292
rect 12880 3236 12936 3292
rect 12936 3236 12940 3292
rect 12876 3232 12940 3236
rect 12956 3292 13020 3296
rect 12956 3236 12960 3292
rect 12960 3236 13016 3292
rect 13016 3236 13020 3292
rect 12956 3232 13020 3236
rect 13036 3292 13100 3296
rect 13036 3236 13040 3292
rect 13040 3236 13096 3292
rect 13096 3236 13100 3292
rect 13036 3232 13100 3236
rect 9260 3224 9324 3228
rect 9260 3168 9310 3224
rect 9310 3168 9324 3224
rect 9260 3164 9324 3168
rect 10548 3028 10612 3092
rect 13492 3028 13556 3092
rect 16068 3028 16132 3092
rect 4108 2756 4172 2820
rect 12388 2756 12452 2820
rect 2926 2748 2990 2752
rect 2926 2692 2930 2748
rect 2930 2692 2986 2748
rect 2986 2692 2990 2748
rect 2926 2688 2990 2692
rect 3006 2748 3070 2752
rect 3006 2692 3010 2748
rect 3010 2692 3066 2748
rect 3066 2692 3070 2748
rect 3006 2688 3070 2692
rect 3086 2748 3150 2752
rect 3086 2692 3090 2748
rect 3090 2692 3146 2748
rect 3146 2692 3150 2748
rect 3086 2688 3150 2692
rect 3166 2748 3230 2752
rect 3166 2692 3170 2748
rect 3170 2692 3226 2748
rect 3226 2692 3230 2748
rect 3166 2688 3230 2692
rect 6874 2748 6938 2752
rect 6874 2692 6878 2748
rect 6878 2692 6934 2748
rect 6934 2692 6938 2748
rect 6874 2688 6938 2692
rect 6954 2748 7018 2752
rect 6954 2692 6958 2748
rect 6958 2692 7014 2748
rect 7014 2692 7018 2748
rect 6954 2688 7018 2692
rect 7034 2748 7098 2752
rect 7034 2692 7038 2748
rect 7038 2692 7094 2748
rect 7094 2692 7098 2748
rect 7034 2688 7098 2692
rect 7114 2748 7178 2752
rect 7114 2692 7118 2748
rect 7118 2692 7174 2748
rect 7174 2692 7178 2748
rect 7114 2688 7178 2692
rect 10822 2748 10886 2752
rect 10822 2692 10826 2748
rect 10826 2692 10882 2748
rect 10882 2692 10886 2748
rect 10822 2688 10886 2692
rect 10902 2748 10966 2752
rect 10902 2692 10906 2748
rect 10906 2692 10962 2748
rect 10962 2692 10966 2748
rect 10902 2688 10966 2692
rect 10982 2748 11046 2752
rect 10982 2692 10986 2748
rect 10986 2692 11042 2748
rect 11042 2692 11046 2748
rect 10982 2688 11046 2692
rect 11062 2748 11126 2752
rect 11062 2692 11066 2748
rect 11066 2692 11122 2748
rect 11122 2692 11126 2748
rect 11062 2688 11126 2692
rect 14770 2748 14834 2752
rect 14770 2692 14774 2748
rect 14774 2692 14830 2748
rect 14830 2692 14834 2748
rect 14770 2688 14834 2692
rect 14850 2748 14914 2752
rect 14850 2692 14854 2748
rect 14854 2692 14910 2748
rect 14910 2692 14914 2748
rect 14850 2688 14914 2692
rect 14930 2748 14994 2752
rect 14930 2692 14934 2748
rect 14934 2692 14990 2748
rect 14990 2692 14994 2748
rect 14930 2688 14994 2692
rect 15010 2748 15074 2752
rect 15010 2692 15014 2748
rect 15014 2692 15070 2748
rect 15070 2692 15074 2748
rect 15010 2688 15074 2692
rect 10180 2620 10244 2684
rect 12204 2620 12268 2684
rect 9812 2484 9876 2548
rect 7788 2212 7852 2276
rect 8156 2212 8220 2276
rect 15332 2348 15396 2412
rect 4900 2204 4964 2208
rect 4900 2148 4904 2204
rect 4904 2148 4960 2204
rect 4960 2148 4964 2204
rect 4900 2144 4964 2148
rect 4980 2204 5044 2208
rect 4980 2148 4984 2204
rect 4984 2148 5040 2204
rect 5040 2148 5044 2204
rect 4980 2144 5044 2148
rect 5060 2204 5124 2208
rect 5060 2148 5064 2204
rect 5064 2148 5120 2204
rect 5120 2148 5124 2204
rect 5060 2144 5124 2148
rect 5140 2204 5204 2208
rect 5140 2148 5144 2204
rect 5144 2148 5200 2204
rect 5200 2148 5204 2204
rect 5140 2144 5204 2148
rect 8848 2204 8912 2208
rect 8848 2148 8852 2204
rect 8852 2148 8908 2204
rect 8908 2148 8912 2204
rect 8848 2144 8912 2148
rect 8928 2204 8992 2208
rect 8928 2148 8932 2204
rect 8932 2148 8988 2204
rect 8988 2148 8992 2204
rect 8928 2144 8992 2148
rect 9008 2204 9072 2208
rect 9008 2148 9012 2204
rect 9012 2148 9068 2204
rect 9068 2148 9072 2204
rect 9008 2144 9072 2148
rect 9088 2204 9152 2208
rect 9088 2148 9092 2204
rect 9092 2148 9148 2204
rect 9148 2148 9152 2204
rect 9088 2144 9152 2148
rect 12796 2204 12860 2208
rect 12796 2148 12800 2204
rect 12800 2148 12856 2204
rect 12856 2148 12860 2204
rect 12796 2144 12860 2148
rect 12876 2204 12940 2208
rect 12876 2148 12880 2204
rect 12880 2148 12936 2204
rect 12936 2148 12940 2204
rect 12876 2144 12940 2148
rect 12956 2204 13020 2208
rect 12956 2148 12960 2204
rect 12960 2148 13016 2204
rect 13016 2148 13020 2204
rect 12956 2144 13020 2148
rect 13036 2204 13100 2208
rect 13036 2148 13040 2204
rect 13040 2148 13096 2204
rect 13096 2148 13100 2204
rect 13036 2144 13100 2148
rect 9444 2076 9508 2140
rect 10364 2076 10428 2140
rect 12388 2136 12452 2140
rect 12388 2080 12438 2136
rect 12438 2080 12452 2136
rect 12388 2076 12452 2080
rect 13676 1804 13740 1868
rect 11468 1668 11532 1732
rect 12572 1668 12636 1732
rect 2926 1660 2990 1664
rect 2926 1604 2930 1660
rect 2930 1604 2986 1660
rect 2986 1604 2990 1660
rect 2926 1600 2990 1604
rect 3006 1660 3070 1664
rect 3006 1604 3010 1660
rect 3010 1604 3066 1660
rect 3066 1604 3070 1660
rect 3006 1600 3070 1604
rect 3086 1660 3150 1664
rect 3086 1604 3090 1660
rect 3090 1604 3146 1660
rect 3146 1604 3150 1660
rect 3086 1600 3150 1604
rect 3166 1660 3230 1664
rect 3166 1604 3170 1660
rect 3170 1604 3226 1660
rect 3226 1604 3230 1660
rect 3166 1600 3230 1604
rect 6874 1660 6938 1664
rect 6874 1604 6878 1660
rect 6878 1604 6934 1660
rect 6934 1604 6938 1660
rect 6874 1600 6938 1604
rect 6954 1660 7018 1664
rect 6954 1604 6958 1660
rect 6958 1604 7014 1660
rect 7014 1604 7018 1660
rect 6954 1600 7018 1604
rect 7034 1660 7098 1664
rect 7034 1604 7038 1660
rect 7038 1604 7094 1660
rect 7094 1604 7098 1660
rect 7034 1600 7098 1604
rect 7114 1660 7178 1664
rect 7114 1604 7118 1660
rect 7118 1604 7174 1660
rect 7174 1604 7178 1660
rect 7114 1600 7178 1604
rect 10822 1660 10886 1664
rect 10822 1604 10826 1660
rect 10826 1604 10882 1660
rect 10882 1604 10886 1660
rect 10822 1600 10886 1604
rect 10902 1660 10966 1664
rect 10902 1604 10906 1660
rect 10906 1604 10962 1660
rect 10962 1604 10966 1660
rect 10902 1600 10966 1604
rect 10982 1660 11046 1664
rect 10982 1604 10986 1660
rect 10986 1604 11042 1660
rect 11042 1604 11046 1660
rect 10982 1600 11046 1604
rect 11062 1660 11126 1664
rect 11062 1604 11066 1660
rect 11066 1604 11122 1660
rect 11122 1604 11126 1660
rect 11062 1600 11126 1604
rect 14770 1660 14834 1664
rect 14770 1604 14774 1660
rect 14774 1604 14830 1660
rect 14830 1604 14834 1660
rect 14770 1600 14834 1604
rect 14850 1660 14914 1664
rect 14850 1604 14854 1660
rect 14854 1604 14910 1660
rect 14910 1604 14914 1660
rect 14850 1600 14914 1604
rect 14930 1660 14994 1664
rect 14930 1604 14934 1660
rect 14934 1604 14990 1660
rect 14990 1604 14994 1660
rect 14930 1600 14994 1604
rect 15010 1660 15074 1664
rect 15010 1604 15014 1660
rect 15014 1604 15070 1660
rect 15070 1604 15074 1660
rect 15010 1600 15074 1604
rect 13492 1532 13556 1596
rect 8156 1396 8220 1460
rect 4900 1116 4964 1120
rect 4900 1060 4904 1116
rect 4904 1060 4960 1116
rect 4960 1060 4964 1116
rect 4900 1056 4964 1060
rect 4980 1116 5044 1120
rect 4980 1060 4984 1116
rect 4984 1060 5040 1116
rect 5040 1060 5044 1116
rect 4980 1056 5044 1060
rect 5060 1116 5124 1120
rect 5060 1060 5064 1116
rect 5064 1060 5120 1116
rect 5120 1060 5124 1116
rect 5060 1056 5124 1060
rect 5140 1116 5204 1120
rect 5140 1060 5144 1116
rect 5144 1060 5200 1116
rect 5200 1060 5204 1116
rect 5140 1056 5204 1060
rect 8848 1116 8912 1120
rect 8848 1060 8852 1116
rect 8852 1060 8908 1116
rect 8908 1060 8912 1116
rect 8848 1056 8912 1060
rect 8928 1116 8992 1120
rect 8928 1060 8932 1116
rect 8932 1060 8988 1116
rect 8988 1060 8992 1116
rect 8928 1056 8992 1060
rect 9008 1116 9072 1120
rect 9008 1060 9012 1116
rect 9012 1060 9068 1116
rect 9068 1060 9072 1116
rect 9008 1056 9072 1060
rect 9088 1116 9152 1120
rect 9088 1060 9092 1116
rect 9092 1060 9148 1116
rect 9148 1060 9152 1116
rect 9088 1056 9152 1060
rect 12796 1116 12860 1120
rect 12796 1060 12800 1116
rect 12800 1060 12856 1116
rect 12856 1060 12860 1116
rect 12796 1056 12860 1060
rect 12876 1116 12940 1120
rect 12876 1060 12880 1116
rect 12880 1060 12936 1116
rect 12936 1060 12940 1116
rect 12876 1056 12940 1060
rect 12956 1116 13020 1120
rect 12956 1060 12960 1116
rect 12960 1060 13016 1116
rect 13016 1060 13020 1116
rect 12956 1056 13020 1060
rect 13036 1116 13100 1120
rect 13036 1060 13040 1116
rect 13040 1060 13096 1116
rect 13096 1060 13100 1116
rect 13036 1056 13100 1060
rect 9444 580 9508 644
rect 13860 580 13924 644
<< metal4 >>
rect 2918 22336 3238 22896
rect 2918 22272 2926 22336
rect 2990 22272 3006 22336
rect 3070 22272 3086 22336
rect 3150 22272 3166 22336
rect 3230 22272 3238 22336
rect 2918 21248 3238 22272
rect 2918 21184 2926 21248
rect 2990 21184 3006 21248
rect 3070 21184 3086 21248
rect 3150 21184 3166 21248
rect 3230 21184 3238 21248
rect 2918 20160 3238 21184
rect 4892 22880 5212 22896
rect 4892 22816 4900 22880
rect 4964 22816 4980 22880
rect 5044 22816 5060 22880
rect 5124 22816 5140 22880
rect 5204 22816 5212 22880
rect 4892 21792 5212 22816
rect 4892 21728 4900 21792
rect 4964 21728 4980 21792
rect 5044 21728 5060 21792
rect 5124 21728 5140 21792
rect 5204 21728 5212 21792
rect 4892 20704 5212 21728
rect 4892 20640 4900 20704
rect 4964 20640 4980 20704
rect 5044 20640 5060 20704
rect 5124 20640 5140 20704
rect 5204 20640 5212 20704
rect 3739 20364 3805 20365
rect 3739 20300 3740 20364
rect 3804 20300 3805 20364
rect 3739 20299 3805 20300
rect 2918 20096 2926 20160
rect 2990 20096 3006 20160
rect 3070 20096 3086 20160
rect 3150 20096 3166 20160
rect 3230 20096 3238 20160
rect 2918 19072 3238 20096
rect 2918 19008 2926 19072
rect 2990 19008 3006 19072
rect 3070 19008 3086 19072
rect 3150 19008 3166 19072
rect 3230 19008 3238 19072
rect 2451 18596 2517 18597
rect 2451 18532 2452 18596
rect 2516 18532 2517 18596
rect 2451 18531 2517 18532
rect 1715 18324 1781 18325
rect 1715 18260 1716 18324
rect 1780 18260 1781 18324
rect 1715 18259 1781 18260
rect 1718 12205 1778 18259
rect 2454 16693 2514 18531
rect 2918 17984 3238 19008
rect 2918 17920 2926 17984
rect 2990 17920 3006 17984
rect 3070 17920 3086 17984
rect 3150 17920 3166 17984
rect 3230 17920 3238 17984
rect 2918 16896 3238 17920
rect 2918 16832 2926 16896
rect 2990 16832 3006 16896
rect 3070 16832 3086 16896
rect 3150 16832 3166 16896
rect 3230 16832 3238 16896
rect 2451 16692 2517 16693
rect 2451 16628 2452 16692
rect 2516 16628 2517 16692
rect 2451 16627 2517 16628
rect 2267 16556 2333 16557
rect 2267 16492 2268 16556
rect 2332 16492 2333 16556
rect 2267 16491 2333 16492
rect 1899 15332 1965 15333
rect 1899 15268 1900 15332
rect 1964 15268 1965 15332
rect 1899 15267 1965 15268
rect 1715 12204 1781 12205
rect 1715 12140 1716 12204
rect 1780 12140 1781 12204
rect 1715 12139 1781 12140
rect 1902 10709 1962 15267
rect 2270 14653 2330 16491
rect 2454 16013 2514 16627
rect 2635 16420 2701 16421
rect 2635 16356 2636 16420
rect 2700 16356 2701 16420
rect 2635 16355 2701 16356
rect 2451 16012 2517 16013
rect 2451 15948 2452 16012
rect 2516 15948 2517 16012
rect 2451 15947 2517 15948
rect 2267 14652 2333 14653
rect 2267 14588 2268 14652
rect 2332 14588 2333 14652
rect 2267 14587 2333 14588
rect 2267 14380 2333 14381
rect 2267 14316 2268 14380
rect 2332 14316 2333 14380
rect 2267 14315 2333 14316
rect 2270 11797 2330 14315
rect 2267 11796 2333 11797
rect 2267 11732 2268 11796
rect 2332 11732 2333 11796
rect 2267 11731 2333 11732
rect 2454 11117 2514 15947
rect 2638 11933 2698 16355
rect 2918 15808 3238 16832
rect 3371 16556 3437 16557
rect 3371 16492 3372 16556
rect 3436 16492 3437 16556
rect 3371 16491 3437 16492
rect 2918 15744 2926 15808
rect 2990 15744 3006 15808
rect 3070 15744 3086 15808
rect 3150 15744 3166 15808
rect 3230 15744 3238 15808
rect 2918 14720 3238 15744
rect 2918 14656 2926 14720
rect 2990 14656 3006 14720
rect 3070 14656 3086 14720
rect 3150 14656 3166 14720
rect 3230 14656 3238 14720
rect 2918 13632 3238 14656
rect 2918 13568 2926 13632
rect 2990 13568 3006 13632
rect 3070 13568 3086 13632
rect 3150 13568 3166 13632
rect 3230 13568 3238 13632
rect 2918 12544 3238 13568
rect 2918 12480 2926 12544
rect 2990 12480 3006 12544
rect 3070 12480 3086 12544
rect 3150 12480 3166 12544
rect 3230 12480 3238 12544
rect 2635 11932 2701 11933
rect 2635 11868 2636 11932
rect 2700 11868 2701 11932
rect 2635 11867 2701 11868
rect 2918 11456 3238 12480
rect 2918 11392 2926 11456
rect 2990 11392 3006 11456
rect 3070 11392 3086 11456
rect 3150 11392 3166 11456
rect 3230 11392 3238 11456
rect 2451 11116 2517 11117
rect 2451 11052 2452 11116
rect 2516 11052 2517 11116
rect 2451 11051 2517 11052
rect 1899 10708 1965 10709
rect 1899 10644 1900 10708
rect 1964 10644 1965 10708
rect 1899 10643 1965 10644
rect 2918 10368 3238 11392
rect 3374 11389 3434 16491
rect 3555 15604 3621 15605
rect 3555 15540 3556 15604
rect 3620 15540 3621 15604
rect 3555 15539 3621 15540
rect 3558 14381 3618 15539
rect 3742 14925 3802 20299
rect 4892 19616 5212 20640
rect 4892 19552 4900 19616
rect 4964 19552 4980 19616
rect 5044 19552 5060 19616
rect 5124 19552 5140 19616
rect 5204 19552 5212 19616
rect 4475 19276 4541 19277
rect 4475 19212 4476 19276
rect 4540 19212 4541 19276
rect 4475 19211 4541 19212
rect 4107 18052 4173 18053
rect 4107 17988 4108 18052
rect 4172 17988 4173 18052
rect 4107 17987 4173 17988
rect 3923 17236 3989 17237
rect 3923 17172 3924 17236
rect 3988 17172 3989 17236
rect 3923 17171 3989 17172
rect 3739 14924 3805 14925
rect 3739 14860 3740 14924
rect 3804 14860 3805 14924
rect 3739 14859 3805 14860
rect 3739 14788 3805 14789
rect 3739 14724 3740 14788
rect 3804 14724 3805 14788
rect 3739 14723 3805 14724
rect 3555 14380 3621 14381
rect 3555 14316 3556 14380
rect 3620 14316 3621 14380
rect 3555 14315 3621 14316
rect 3555 14244 3621 14245
rect 3555 14180 3556 14244
rect 3620 14180 3621 14244
rect 3555 14179 3621 14180
rect 3558 12885 3618 14179
rect 3742 13021 3802 14723
rect 3926 14381 3986 17171
rect 3923 14380 3989 14381
rect 3923 14316 3924 14380
rect 3988 14316 3989 14380
rect 3923 14315 3989 14316
rect 3739 13020 3805 13021
rect 3739 12956 3740 13020
rect 3804 12956 3805 13020
rect 3739 12955 3805 12956
rect 3555 12884 3621 12885
rect 3555 12820 3556 12884
rect 3620 12820 3621 12884
rect 3555 12819 3621 12820
rect 3923 12884 3989 12885
rect 3923 12820 3924 12884
rect 3988 12820 3989 12884
rect 3923 12819 3989 12820
rect 3555 12612 3621 12613
rect 3555 12548 3556 12612
rect 3620 12548 3621 12612
rect 3555 12547 3621 12548
rect 3739 12612 3805 12613
rect 3739 12548 3740 12612
rect 3804 12548 3805 12612
rect 3739 12547 3805 12548
rect 3371 11388 3437 11389
rect 3371 11324 3372 11388
rect 3436 11324 3437 11388
rect 3371 11323 3437 11324
rect 3558 11253 3618 12547
rect 3742 12205 3802 12547
rect 3739 12204 3805 12205
rect 3739 12140 3740 12204
rect 3804 12140 3805 12204
rect 3739 12139 3805 12140
rect 3739 12068 3805 12069
rect 3739 12004 3740 12068
rect 3804 12004 3805 12068
rect 3739 12003 3805 12004
rect 3555 11252 3621 11253
rect 3555 11188 3556 11252
rect 3620 11188 3621 11252
rect 3555 11187 3621 11188
rect 2918 10304 2926 10368
rect 2990 10304 3006 10368
rect 3070 10304 3086 10368
rect 3150 10304 3166 10368
rect 3230 10304 3238 10368
rect 2918 9280 3238 10304
rect 3742 9485 3802 12003
rect 3926 10981 3986 12819
rect 3923 10980 3989 10981
rect 3923 10916 3924 10980
rect 3988 10916 3989 10980
rect 3923 10915 3989 10916
rect 4110 10437 4170 17987
rect 4291 15876 4357 15877
rect 4291 15812 4292 15876
rect 4356 15812 4357 15876
rect 4291 15811 4357 15812
rect 4294 12477 4354 15811
rect 4478 14925 4538 19211
rect 4659 18868 4725 18869
rect 4659 18804 4660 18868
rect 4724 18804 4725 18868
rect 4659 18803 4725 18804
rect 4475 14924 4541 14925
rect 4475 14860 4476 14924
rect 4540 14860 4541 14924
rect 4475 14859 4541 14860
rect 4475 14652 4541 14653
rect 4475 14588 4476 14652
rect 4540 14588 4541 14652
rect 4475 14587 4541 14588
rect 4478 13701 4538 14587
rect 4475 13700 4541 13701
rect 4475 13636 4476 13700
rect 4540 13636 4541 13700
rect 4475 13635 4541 13636
rect 4475 13428 4541 13429
rect 4475 13364 4476 13428
rect 4540 13364 4541 13428
rect 4475 13363 4541 13364
rect 4291 12476 4357 12477
rect 4291 12412 4292 12476
rect 4356 12412 4357 12476
rect 4291 12411 4357 12412
rect 4291 12340 4357 12341
rect 4291 12276 4292 12340
rect 4356 12276 4357 12340
rect 4291 12275 4357 12276
rect 4294 12069 4354 12275
rect 4291 12068 4357 12069
rect 4291 12004 4292 12068
rect 4356 12004 4357 12068
rect 4291 12003 4357 12004
rect 4291 11932 4357 11933
rect 4291 11868 4292 11932
rect 4356 11868 4357 11932
rect 4291 11867 4357 11868
rect 4107 10436 4173 10437
rect 4107 10372 4108 10436
rect 4172 10372 4173 10436
rect 4107 10371 4173 10372
rect 4294 10165 4354 11867
rect 4291 10164 4357 10165
rect 4291 10100 4292 10164
rect 4356 10100 4357 10164
rect 4291 10099 4357 10100
rect 3739 9484 3805 9485
rect 3739 9420 3740 9484
rect 3804 9420 3805 9484
rect 3739 9419 3805 9420
rect 2918 9216 2926 9280
rect 2990 9216 3006 9280
rect 3070 9216 3086 9280
rect 3150 9216 3166 9280
rect 3230 9216 3238 9280
rect 2918 8192 3238 9216
rect 4478 8397 4538 13363
rect 4662 13021 4722 18803
rect 4892 18528 5212 19552
rect 6866 22336 7186 22896
rect 6866 22272 6874 22336
rect 6938 22272 6954 22336
rect 7018 22272 7034 22336
rect 7098 22272 7114 22336
rect 7178 22272 7186 22336
rect 6866 21248 7186 22272
rect 6866 21184 6874 21248
rect 6938 21184 6954 21248
rect 7018 21184 7034 21248
rect 7098 21184 7114 21248
rect 7178 21184 7186 21248
rect 6866 20160 7186 21184
rect 6866 20096 6874 20160
rect 6938 20096 6954 20160
rect 7018 20096 7034 20160
rect 7098 20096 7114 20160
rect 7178 20096 7186 20160
rect 6866 19072 7186 20096
rect 6866 19008 6874 19072
rect 6938 19008 6954 19072
rect 7018 19008 7034 19072
rect 7098 19008 7114 19072
rect 7178 19008 7186 19072
rect 5763 18732 5829 18733
rect 5763 18668 5764 18732
rect 5828 18668 5829 18732
rect 5763 18667 5829 18668
rect 4892 18464 4900 18528
rect 4964 18464 4980 18528
rect 5044 18464 5060 18528
rect 5124 18464 5140 18528
rect 5204 18464 5212 18528
rect 4892 17440 5212 18464
rect 4892 17376 4900 17440
rect 4964 17376 4980 17440
rect 5044 17376 5060 17440
rect 5124 17376 5140 17440
rect 5204 17376 5212 17440
rect 4892 16352 5212 17376
rect 5395 16828 5461 16829
rect 5395 16764 5396 16828
rect 5460 16764 5461 16828
rect 5395 16763 5461 16764
rect 4892 16288 4900 16352
rect 4964 16288 4980 16352
rect 5044 16288 5060 16352
rect 5124 16288 5140 16352
rect 5204 16288 5212 16352
rect 4892 15264 5212 16288
rect 5398 15877 5458 16763
rect 5579 16556 5645 16557
rect 5579 16492 5580 16556
rect 5644 16492 5645 16556
rect 5579 16491 5645 16492
rect 5395 15876 5461 15877
rect 5395 15812 5396 15876
rect 5460 15812 5461 15876
rect 5395 15811 5461 15812
rect 5395 15332 5461 15333
rect 5395 15268 5396 15332
rect 5460 15268 5461 15332
rect 5395 15267 5461 15268
rect 4892 15200 4900 15264
rect 4964 15200 4980 15264
rect 5044 15200 5060 15264
rect 5124 15200 5140 15264
rect 5204 15200 5212 15264
rect 4892 14176 5212 15200
rect 4892 14112 4900 14176
rect 4964 14112 4980 14176
rect 5044 14112 5060 14176
rect 5124 14112 5140 14176
rect 5204 14112 5212 14176
rect 4892 13088 5212 14112
rect 4892 13024 4900 13088
rect 4964 13024 4980 13088
rect 5044 13024 5060 13088
rect 5124 13024 5140 13088
rect 5204 13024 5212 13088
rect 4659 13020 4725 13021
rect 4659 12956 4660 13020
rect 4724 12956 4725 13020
rect 4659 12955 4725 12956
rect 4659 12748 4725 12749
rect 4659 12684 4660 12748
rect 4724 12684 4725 12748
rect 4659 12683 4725 12684
rect 4662 11389 4722 12683
rect 4892 12000 5212 13024
rect 4892 11936 4900 12000
rect 4964 11936 4980 12000
rect 5044 11936 5060 12000
rect 5124 11936 5140 12000
rect 5204 11936 5212 12000
rect 4659 11388 4725 11389
rect 4659 11324 4660 11388
rect 4724 11324 4725 11388
rect 4659 11323 4725 11324
rect 4659 10980 4725 10981
rect 4659 10916 4660 10980
rect 4724 10916 4725 10980
rect 4659 10915 4725 10916
rect 4662 8397 4722 10915
rect 4892 10912 5212 11936
rect 5398 11797 5458 15267
rect 5582 13701 5642 16491
rect 5579 13700 5645 13701
rect 5579 13636 5580 13700
rect 5644 13636 5645 13700
rect 5579 13635 5645 13636
rect 5579 13564 5645 13565
rect 5579 13500 5580 13564
rect 5644 13500 5645 13564
rect 5579 13499 5645 13500
rect 5395 11796 5461 11797
rect 5395 11732 5396 11796
rect 5460 11732 5461 11796
rect 5395 11731 5461 11732
rect 4892 10848 4900 10912
rect 4964 10848 4980 10912
rect 5044 10848 5060 10912
rect 5124 10848 5140 10912
rect 5204 10848 5212 10912
rect 4892 9824 5212 10848
rect 5582 10573 5642 13499
rect 5766 12749 5826 18667
rect 5947 18324 6013 18325
rect 5947 18260 5948 18324
rect 6012 18260 6013 18324
rect 5947 18259 6013 18260
rect 5950 14109 6010 18259
rect 6131 18052 6197 18053
rect 6131 17988 6132 18052
rect 6196 17988 6197 18052
rect 6131 17987 6197 17988
rect 6134 15197 6194 17987
rect 6866 17984 7186 19008
rect 8840 22880 9160 22896
rect 8840 22816 8848 22880
rect 8912 22816 8928 22880
rect 8992 22816 9008 22880
rect 9072 22816 9088 22880
rect 9152 22816 9160 22880
rect 8840 21792 9160 22816
rect 8840 21728 8848 21792
rect 8912 21728 8928 21792
rect 8992 21728 9008 21792
rect 9072 21728 9088 21792
rect 9152 21728 9160 21792
rect 8840 20704 9160 21728
rect 8840 20640 8848 20704
rect 8912 20640 8928 20704
rect 8992 20640 9008 20704
rect 9072 20640 9088 20704
rect 9152 20640 9160 20704
rect 8840 19616 9160 20640
rect 8840 19552 8848 19616
rect 8912 19552 8928 19616
rect 8992 19552 9008 19616
rect 9072 19552 9088 19616
rect 9152 19552 9160 19616
rect 8840 18528 9160 19552
rect 8840 18464 8848 18528
rect 8912 18464 8928 18528
rect 8992 18464 9008 18528
rect 9072 18464 9088 18528
rect 9152 18464 9160 18528
rect 8707 18460 8773 18461
rect 8707 18396 8708 18460
rect 8772 18396 8773 18460
rect 8707 18395 8773 18396
rect 7787 18324 7853 18325
rect 7787 18260 7788 18324
rect 7852 18260 7853 18324
rect 7787 18259 7853 18260
rect 6866 17920 6874 17984
rect 6938 17920 6954 17984
rect 7018 17920 7034 17984
rect 7098 17920 7114 17984
rect 7178 17920 7186 17984
rect 6499 17100 6565 17101
rect 6499 17036 6500 17100
rect 6564 17036 6565 17100
rect 6499 17035 6565 17036
rect 6315 16284 6381 16285
rect 6315 16220 6316 16284
rect 6380 16220 6381 16284
rect 6315 16219 6381 16220
rect 6131 15196 6197 15197
rect 6131 15132 6132 15196
rect 6196 15132 6197 15196
rect 6131 15131 6197 15132
rect 6131 15060 6197 15061
rect 6131 14996 6132 15060
rect 6196 14996 6197 15060
rect 6131 14995 6197 14996
rect 5947 14108 6013 14109
rect 5947 14044 5948 14108
rect 6012 14044 6013 14108
rect 5947 14043 6013 14044
rect 5950 13157 6010 14043
rect 5947 13156 6013 13157
rect 5947 13092 5948 13156
rect 6012 13092 6013 13156
rect 5947 13091 6013 13092
rect 6134 13018 6194 14995
rect 5950 12958 6194 13018
rect 5763 12748 5829 12749
rect 5763 12684 5764 12748
rect 5828 12684 5829 12748
rect 5763 12683 5829 12684
rect 5950 11253 6010 12958
rect 6131 12884 6197 12885
rect 6131 12820 6132 12884
rect 6196 12820 6197 12884
rect 6131 12819 6197 12820
rect 5947 11252 6013 11253
rect 5947 11188 5948 11252
rect 6012 11188 6013 11252
rect 5947 11187 6013 11188
rect 6134 10573 6194 12819
rect 6318 11525 6378 16219
rect 6502 12477 6562 17035
rect 6866 16896 7186 17920
rect 6866 16832 6874 16896
rect 6938 16832 6954 16896
rect 7018 16832 7034 16896
rect 7098 16832 7114 16896
rect 7178 16832 7186 16896
rect 6683 16420 6749 16421
rect 6683 16356 6684 16420
rect 6748 16356 6749 16420
rect 6683 16355 6749 16356
rect 6499 12476 6565 12477
rect 6499 12412 6500 12476
rect 6564 12412 6565 12476
rect 6499 12411 6565 12412
rect 6686 12205 6746 16355
rect 6866 15808 7186 16832
rect 7603 16692 7669 16693
rect 7603 16628 7604 16692
rect 7668 16628 7669 16692
rect 7603 16627 7669 16628
rect 7419 16556 7485 16557
rect 7419 16492 7420 16556
rect 7484 16492 7485 16556
rect 7419 16491 7485 16492
rect 6866 15744 6874 15808
rect 6938 15744 6954 15808
rect 7018 15744 7034 15808
rect 7098 15744 7114 15808
rect 7178 15744 7186 15808
rect 6866 14720 7186 15744
rect 7281 15740 7347 15741
rect 7281 15676 7282 15740
rect 7346 15676 7347 15740
rect 7281 15675 7347 15676
rect 6866 14656 6874 14720
rect 6938 14656 6954 14720
rect 7018 14656 7034 14720
rect 7098 14656 7114 14720
rect 7178 14656 7186 14720
rect 6866 13632 7186 14656
rect 6866 13568 6874 13632
rect 6938 13568 6954 13632
rect 7018 13568 7034 13632
rect 7098 13568 7114 13632
rect 7178 13568 7186 13632
rect 6866 12544 7186 13568
rect 6866 12480 6874 12544
rect 6938 12480 6954 12544
rect 7018 12480 7034 12544
rect 7098 12480 7114 12544
rect 7178 12480 7186 12544
rect 6683 12204 6749 12205
rect 6683 12140 6684 12204
rect 6748 12140 6749 12204
rect 6683 12139 6749 12140
rect 6315 11524 6381 11525
rect 6315 11460 6316 11524
rect 6380 11460 6381 11524
rect 6315 11459 6381 11460
rect 6866 11456 7186 12480
rect 7284 11933 7344 15675
rect 7281 11932 7347 11933
rect 7281 11868 7282 11932
rect 7346 11868 7347 11932
rect 7281 11867 7347 11868
rect 6866 11392 6874 11456
rect 6938 11392 6954 11456
rect 7018 11392 7034 11456
rect 7098 11392 7114 11456
rect 7178 11392 7186 11456
rect 5579 10572 5645 10573
rect 5579 10508 5580 10572
rect 5644 10508 5645 10572
rect 5579 10507 5645 10508
rect 6131 10572 6197 10573
rect 6131 10508 6132 10572
rect 6196 10508 6197 10572
rect 6131 10507 6197 10508
rect 6866 10368 7186 11392
rect 6866 10304 6874 10368
rect 6938 10304 6954 10368
rect 7018 10304 7034 10368
rect 7098 10304 7114 10368
rect 7178 10304 7186 10368
rect 6131 9892 6197 9893
rect 6131 9828 6132 9892
rect 6196 9828 6197 9892
rect 6131 9827 6197 9828
rect 4892 9760 4900 9824
rect 4964 9760 4980 9824
rect 5044 9760 5060 9824
rect 5124 9760 5140 9824
rect 5204 9760 5212 9824
rect 4892 8736 5212 9760
rect 4892 8672 4900 8736
rect 4964 8672 4980 8736
rect 5044 8672 5060 8736
rect 5124 8672 5140 8736
rect 5204 8672 5212 8736
rect 4475 8396 4541 8397
rect 4475 8332 4476 8396
rect 4540 8332 4541 8396
rect 4475 8331 4541 8332
rect 4659 8396 4725 8397
rect 4659 8332 4660 8396
rect 4724 8332 4725 8396
rect 4659 8331 4725 8332
rect 2918 8128 2926 8192
rect 2990 8128 3006 8192
rect 3070 8128 3086 8192
rect 3150 8128 3166 8192
rect 3230 8128 3238 8192
rect 2918 7104 3238 8128
rect 4291 7852 4357 7853
rect 4291 7788 4292 7852
rect 4356 7788 4357 7852
rect 4291 7787 4357 7788
rect 4107 7444 4173 7445
rect 4107 7380 4108 7444
rect 4172 7380 4173 7444
rect 4107 7379 4173 7380
rect 2918 7040 2926 7104
rect 2990 7040 3006 7104
rect 3070 7040 3086 7104
rect 3150 7040 3166 7104
rect 3230 7040 3238 7104
rect 2635 6900 2701 6901
rect 2635 6836 2636 6900
rect 2700 6836 2701 6900
rect 2635 6835 2701 6836
rect 2638 3501 2698 6835
rect 2918 6016 3238 7040
rect 2918 5952 2926 6016
rect 2990 5952 3006 6016
rect 3070 5952 3086 6016
rect 3150 5952 3166 6016
rect 3230 5952 3238 6016
rect 2918 4928 3238 5952
rect 4110 5677 4170 7379
rect 4107 5676 4173 5677
rect 4107 5612 4108 5676
rect 4172 5612 4173 5676
rect 4107 5611 4173 5612
rect 2918 4864 2926 4928
rect 2990 4864 3006 4928
rect 3070 4864 3086 4928
rect 3150 4864 3166 4928
rect 3230 4864 3238 4928
rect 2918 3840 3238 4864
rect 2918 3776 2926 3840
rect 2990 3776 3006 3840
rect 3070 3776 3086 3840
rect 3150 3776 3166 3840
rect 3230 3776 3238 3840
rect 2635 3500 2701 3501
rect 2635 3436 2636 3500
rect 2700 3436 2701 3500
rect 2635 3435 2701 3436
rect 2918 2752 3238 3776
rect 4110 2821 4170 5611
rect 4294 3365 4354 7787
rect 4892 7648 5212 8672
rect 5763 7988 5829 7989
rect 5763 7924 5764 7988
rect 5828 7924 5829 7988
rect 5763 7923 5829 7924
rect 5579 7716 5645 7717
rect 5579 7652 5580 7716
rect 5644 7652 5645 7716
rect 5579 7651 5645 7652
rect 4892 7584 4900 7648
rect 4964 7584 4980 7648
rect 5044 7584 5060 7648
rect 5124 7584 5140 7648
rect 5204 7584 5212 7648
rect 4892 6560 5212 7584
rect 4892 6496 4900 6560
rect 4964 6496 4980 6560
rect 5044 6496 5060 6560
rect 5124 6496 5140 6560
rect 5204 6496 5212 6560
rect 4892 5472 5212 6496
rect 4892 5408 4900 5472
rect 4964 5408 4980 5472
rect 5044 5408 5060 5472
rect 5124 5408 5140 5472
rect 5204 5408 5212 5472
rect 4892 4384 5212 5408
rect 4892 4320 4900 4384
rect 4964 4320 4980 4384
rect 5044 4320 5060 4384
rect 5124 4320 5140 4384
rect 5204 4320 5212 4384
rect 4291 3364 4357 3365
rect 4291 3300 4292 3364
rect 4356 3300 4357 3364
rect 4291 3299 4357 3300
rect 4892 3296 5212 4320
rect 4892 3232 4900 3296
rect 4964 3232 4980 3296
rect 5044 3232 5060 3296
rect 5124 3232 5140 3296
rect 5204 3232 5212 3296
rect 4107 2820 4173 2821
rect 4107 2756 4108 2820
rect 4172 2756 4173 2820
rect 4107 2755 4173 2756
rect 2918 2688 2926 2752
rect 2990 2688 3006 2752
rect 3070 2688 3086 2752
rect 3150 2688 3166 2752
rect 3230 2688 3238 2752
rect 2918 1664 3238 2688
rect 2918 1600 2926 1664
rect 2990 1600 3006 1664
rect 3070 1600 3086 1664
rect 3150 1600 3166 1664
rect 3230 1600 3238 1664
rect 2918 1040 3238 1600
rect 4892 2208 5212 3232
rect 5582 3229 5642 7651
rect 5766 3773 5826 7923
rect 6134 5133 6194 9827
rect 6683 9348 6749 9349
rect 6683 9284 6684 9348
rect 6748 9284 6749 9348
rect 6683 9283 6749 9284
rect 6315 5812 6381 5813
rect 6315 5748 6316 5812
rect 6380 5748 6381 5812
rect 6315 5747 6381 5748
rect 6131 5132 6197 5133
rect 6131 5068 6132 5132
rect 6196 5068 6197 5132
rect 6131 5067 6197 5068
rect 6318 3909 6378 5747
rect 6686 5269 6746 9283
rect 6866 9280 7186 10304
rect 6866 9216 6874 9280
rect 6938 9216 6954 9280
rect 7018 9216 7034 9280
rect 7098 9216 7114 9280
rect 7178 9216 7186 9280
rect 6866 8192 7186 9216
rect 6866 8128 6874 8192
rect 6938 8128 6954 8192
rect 7018 8128 7034 8192
rect 7098 8128 7114 8192
rect 7178 8128 7186 8192
rect 6866 7104 7186 8128
rect 6866 7040 6874 7104
rect 6938 7040 6954 7104
rect 7018 7040 7034 7104
rect 7098 7040 7114 7104
rect 7178 7040 7186 7104
rect 6866 6016 7186 7040
rect 6866 5952 6874 6016
rect 6938 5952 6954 6016
rect 7018 5952 7034 6016
rect 7098 5952 7114 6016
rect 7178 5952 7186 6016
rect 6683 5268 6749 5269
rect 6683 5204 6684 5268
rect 6748 5204 6749 5268
rect 6683 5203 6749 5204
rect 6866 4928 7186 5952
rect 6866 4864 6874 4928
rect 6938 4864 6954 4928
rect 7018 4864 7034 4928
rect 7098 4864 7114 4928
rect 7178 4864 7186 4928
rect 6315 3908 6381 3909
rect 6315 3844 6316 3908
rect 6380 3844 6381 3908
rect 6315 3843 6381 3844
rect 6866 3840 7186 4864
rect 7422 3909 7482 16491
rect 7606 15333 7666 16627
rect 7603 15332 7669 15333
rect 7603 15268 7604 15332
rect 7668 15268 7669 15332
rect 7603 15267 7669 15268
rect 7606 9757 7666 15267
rect 7790 13565 7850 18259
rect 8155 17916 8221 17917
rect 8155 17852 8156 17916
rect 8220 17852 8221 17916
rect 8155 17851 8221 17852
rect 7971 16964 8037 16965
rect 7971 16900 7972 16964
rect 8036 16900 8037 16964
rect 7971 16899 8037 16900
rect 7974 15741 8034 16899
rect 7971 15740 8037 15741
rect 7971 15676 7972 15740
rect 8036 15676 8037 15740
rect 7971 15675 8037 15676
rect 7971 14788 8037 14789
rect 7971 14724 7972 14788
rect 8036 14724 8037 14788
rect 7971 14723 8037 14724
rect 7787 13564 7853 13565
rect 7787 13500 7788 13564
rect 7852 13500 7853 13564
rect 7787 13499 7853 13500
rect 7790 12613 7850 13499
rect 7787 12612 7853 12613
rect 7787 12548 7788 12612
rect 7852 12548 7853 12612
rect 7787 12547 7853 12548
rect 7974 12338 8034 14723
rect 8158 13021 8218 17851
rect 8710 16829 8770 18395
rect 8840 17440 9160 18464
rect 10814 22336 11134 22896
rect 10814 22272 10822 22336
rect 10886 22272 10902 22336
rect 10966 22272 10982 22336
rect 11046 22272 11062 22336
rect 11126 22272 11134 22336
rect 10814 21248 11134 22272
rect 10814 21184 10822 21248
rect 10886 21184 10902 21248
rect 10966 21184 10982 21248
rect 11046 21184 11062 21248
rect 11126 21184 11134 21248
rect 10814 20160 11134 21184
rect 10814 20096 10822 20160
rect 10886 20096 10902 20160
rect 10966 20096 10982 20160
rect 11046 20096 11062 20160
rect 11126 20096 11134 20160
rect 10814 19072 11134 20096
rect 10814 19008 10822 19072
rect 10886 19008 10902 19072
rect 10966 19008 10982 19072
rect 11046 19008 11062 19072
rect 11126 19008 11134 19072
rect 9259 18052 9325 18053
rect 9259 17988 9260 18052
rect 9324 17988 9325 18052
rect 9259 17987 9325 17988
rect 9811 18052 9877 18053
rect 9811 17988 9812 18052
rect 9876 17988 9877 18052
rect 9811 17987 9877 17988
rect 8840 17376 8848 17440
rect 8912 17376 8928 17440
rect 8992 17376 9008 17440
rect 9072 17376 9088 17440
rect 9152 17376 9160 17440
rect 8707 16828 8773 16829
rect 8707 16764 8708 16828
rect 8772 16764 8773 16828
rect 8707 16763 8773 16764
rect 8523 16692 8589 16693
rect 8523 16628 8524 16692
rect 8588 16628 8589 16692
rect 8523 16627 8589 16628
rect 8339 15604 8405 15605
rect 8339 15540 8340 15604
rect 8404 15540 8405 15604
rect 8339 15539 8405 15540
rect 8155 13020 8221 13021
rect 8155 12956 8156 13020
rect 8220 12956 8221 13020
rect 8155 12955 8221 12956
rect 8155 12612 8221 12613
rect 8155 12548 8156 12612
rect 8220 12548 8221 12612
rect 8155 12547 8221 12548
rect 7790 12278 8034 12338
rect 7790 10573 7850 12278
rect 7971 12204 8037 12205
rect 7971 12140 7972 12204
rect 8036 12140 8037 12204
rect 7971 12139 8037 12140
rect 7787 10572 7853 10573
rect 7787 10508 7788 10572
rect 7852 10508 7853 10572
rect 7787 10507 7853 10508
rect 7603 9756 7669 9757
rect 7603 9692 7604 9756
rect 7668 9692 7669 9756
rect 7603 9691 7669 9692
rect 7603 8124 7669 8125
rect 7603 8060 7604 8124
rect 7668 8060 7669 8124
rect 7603 8059 7669 8060
rect 7419 3908 7485 3909
rect 7419 3844 7420 3908
rect 7484 3844 7485 3908
rect 7419 3843 7485 3844
rect 6866 3776 6874 3840
rect 6938 3776 6954 3840
rect 7018 3776 7034 3840
rect 7098 3776 7114 3840
rect 7178 3776 7186 3840
rect 5763 3772 5829 3773
rect 5763 3708 5764 3772
rect 5828 3708 5829 3772
rect 5763 3707 5829 3708
rect 5579 3228 5645 3229
rect 5579 3164 5580 3228
rect 5644 3164 5645 3228
rect 5579 3163 5645 3164
rect 4892 2144 4900 2208
rect 4964 2144 4980 2208
rect 5044 2144 5060 2208
rect 5124 2144 5140 2208
rect 5204 2144 5212 2208
rect 4892 1120 5212 2144
rect 4892 1056 4900 1120
rect 4964 1056 4980 1120
rect 5044 1056 5060 1120
rect 5124 1056 5140 1120
rect 5204 1056 5212 1120
rect 4892 1040 5212 1056
rect 6866 2752 7186 3776
rect 7606 3365 7666 8059
rect 7790 4589 7850 10507
rect 7974 5405 8034 12139
rect 8158 11525 8218 12547
rect 8155 11524 8221 11525
rect 8155 11460 8156 11524
rect 8220 11460 8221 11524
rect 8155 11459 8221 11460
rect 8155 11252 8221 11253
rect 8155 11188 8156 11252
rect 8220 11188 8221 11252
rect 8155 11187 8221 11188
rect 8158 8261 8218 11187
rect 8155 8260 8221 8261
rect 8155 8196 8156 8260
rect 8220 8196 8221 8260
rect 8155 8195 8221 8196
rect 8155 6492 8221 6493
rect 8155 6428 8156 6492
rect 8220 6428 8221 6492
rect 8155 6427 8221 6428
rect 7971 5404 8037 5405
rect 7971 5340 7972 5404
rect 8036 5340 8037 5404
rect 7971 5339 8037 5340
rect 7787 4588 7853 4589
rect 7787 4524 7788 4588
rect 7852 4524 7853 4588
rect 7787 4523 7853 4524
rect 7971 4180 8037 4181
rect 7971 4116 7972 4180
rect 8036 4116 8037 4180
rect 7971 4115 8037 4116
rect 7787 3908 7853 3909
rect 7787 3844 7788 3908
rect 7852 3844 7853 3908
rect 7787 3843 7853 3844
rect 7603 3364 7669 3365
rect 7603 3300 7604 3364
rect 7668 3300 7669 3364
rect 7603 3299 7669 3300
rect 6866 2688 6874 2752
rect 6938 2688 6954 2752
rect 7018 2688 7034 2752
rect 7098 2688 7114 2752
rect 7178 2688 7186 2752
rect 6866 1664 7186 2688
rect 7790 2277 7850 3843
rect 7974 3501 8034 4115
rect 7971 3500 8037 3501
rect 7971 3436 7972 3500
rect 8036 3436 8037 3500
rect 7971 3435 8037 3436
rect 8158 2277 8218 6427
rect 8342 3773 8402 15539
rect 8526 11661 8586 16627
rect 8840 16352 9160 17376
rect 8840 16288 8848 16352
rect 8912 16288 8928 16352
rect 8992 16288 9008 16352
rect 9072 16288 9088 16352
rect 9152 16288 9160 16352
rect 8707 15876 8773 15877
rect 8707 15812 8708 15876
rect 8772 15812 8773 15876
rect 8707 15811 8773 15812
rect 8710 13837 8770 15811
rect 8840 15264 9160 16288
rect 8840 15200 8848 15264
rect 8912 15200 8928 15264
rect 8992 15200 9008 15264
rect 9072 15200 9088 15264
rect 9152 15200 9160 15264
rect 8840 14176 9160 15200
rect 9262 14789 9322 17987
rect 9814 17101 9874 17987
rect 10814 17984 11134 19008
rect 12788 22880 13108 22896
rect 12788 22816 12796 22880
rect 12860 22816 12876 22880
rect 12940 22816 12956 22880
rect 13020 22816 13036 22880
rect 13100 22816 13108 22880
rect 12788 21792 13108 22816
rect 12788 21728 12796 21792
rect 12860 21728 12876 21792
rect 12940 21728 12956 21792
rect 13020 21728 13036 21792
rect 13100 21728 13108 21792
rect 12788 20704 13108 21728
rect 12788 20640 12796 20704
rect 12860 20640 12876 20704
rect 12940 20640 12956 20704
rect 13020 20640 13036 20704
rect 13100 20640 13108 20704
rect 12788 19616 13108 20640
rect 12788 19552 12796 19616
rect 12860 19552 12876 19616
rect 12940 19552 12956 19616
rect 13020 19552 13036 19616
rect 13100 19552 13108 19616
rect 12788 18528 13108 19552
rect 12788 18464 12796 18528
rect 12860 18464 12876 18528
rect 12940 18464 12956 18528
rect 13020 18464 13036 18528
rect 13100 18464 13108 18528
rect 11467 18460 11533 18461
rect 11467 18396 11468 18460
rect 11532 18396 11533 18460
rect 11467 18395 11533 18396
rect 10814 17920 10822 17984
rect 10886 17920 10902 17984
rect 10966 17920 10982 17984
rect 11046 17920 11062 17984
rect 11126 17920 11134 17984
rect 10547 17372 10613 17373
rect 10547 17308 10548 17372
rect 10612 17308 10613 17372
rect 10547 17307 10613 17308
rect 9443 17100 9509 17101
rect 9443 17036 9444 17100
rect 9508 17036 9509 17100
rect 9443 17035 9509 17036
rect 9811 17100 9877 17101
rect 9811 17036 9812 17100
rect 9876 17036 9877 17100
rect 9811 17035 9877 17036
rect 9259 14788 9325 14789
rect 9259 14724 9260 14788
rect 9324 14724 9325 14788
rect 9259 14723 9325 14724
rect 8840 14112 8848 14176
rect 8912 14112 8928 14176
rect 8992 14112 9008 14176
rect 9072 14112 9088 14176
rect 9152 14112 9160 14176
rect 8707 13836 8773 13837
rect 8707 13772 8708 13836
rect 8772 13772 8773 13836
rect 8707 13771 8773 13772
rect 8707 13564 8773 13565
rect 8707 13500 8708 13564
rect 8772 13500 8773 13564
rect 8707 13499 8773 13500
rect 8710 12477 8770 13499
rect 8840 13088 9160 14112
rect 8840 13024 8848 13088
rect 8912 13024 8928 13088
rect 8992 13024 9008 13088
rect 9072 13024 9088 13088
rect 9152 13024 9160 13088
rect 8707 12476 8773 12477
rect 8707 12412 8708 12476
rect 8772 12412 8773 12476
rect 8707 12411 8773 12412
rect 8707 12068 8773 12069
rect 8707 12004 8708 12068
rect 8772 12004 8773 12068
rect 8707 12003 8773 12004
rect 8710 11661 8770 12003
rect 8840 12000 9160 13024
rect 8840 11936 8848 12000
rect 8912 11936 8928 12000
rect 8992 11936 9008 12000
rect 9072 11936 9088 12000
rect 9152 11936 9160 12000
rect 8523 11660 8589 11661
rect 8523 11596 8524 11660
rect 8588 11596 8589 11660
rect 8523 11595 8589 11596
rect 8707 11660 8773 11661
rect 8707 11596 8708 11660
rect 8772 11596 8773 11660
rect 8707 11595 8773 11596
rect 8523 11524 8589 11525
rect 8523 11460 8524 11524
rect 8588 11460 8589 11524
rect 8523 11459 8589 11460
rect 8526 10165 8586 11459
rect 8707 10980 8773 10981
rect 8707 10916 8708 10980
rect 8772 10916 8773 10980
rect 8707 10915 8773 10916
rect 8523 10164 8589 10165
rect 8523 10100 8524 10164
rect 8588 10100 8589 10164
rect 8523 10099 8589 10100
rect 8526 6357 8586 10099
rect 8523 6356 8589 6357
rect 8523 6292 8524 6356
rect 8588 6292 8589 6356
rect 8523 6291 8589 6292
rect 8339 3772 8405 3773
rect 8339 3708 8340 3772
rect 8404 3708 8405 3772
rect 8339 3707 8405 3708
rect 8526 3365 8586 6291
rect 8710 4861 8770 10915
rect 8840 10912 9160 11936
rect 9262 11389 9322 14723
rect 9446 12749 9506 17035
rect 9811 16420 9877 16421
rect 9811 16356 9812 16420
rect 9876 16356 9877 16420
rect 9811 16355 9877 16356
rect 9995 16420 10061 16421
rect 9995 16356 9996 16420
rect 10060 16356 10061 16420
rect 9995 16355 10061 16356
rect 9814 15469 9874 16355
rect 9811 15468 9877 15469
rect 9811 15404 9812 15468
rect 9876 15404 9877 15468
rect 9811 15403 9877 15404
rect 9811 15060 9877 15061
rect 9811 14996 9812 15060
rect 9876 14996 9877 15060
rect 9811 14995 9877 14996
rect 9627 14380 9693 14381
rect 9627 14316 9628 14380
rect 9692 14316 9693 14380
rect 9627 14315 9693 14316
rect 9443 12748 9509 12749
rect 9443 12684 9444 12748
rect 9508 12684 9509 12748
rect 9443 12683 9509 12684
rect 9443 12612 9509 12613
rect 9443 12548 9444 12612
rect 9508 12548 9509 12612
rect 9443 12547 9509 12548
rect 9259 11388 9325 11389
rect 9259 11324 9260 11388
rect 9324 11324 9325 11388
rect 9259 11323 9325 11324
rect 8840 10848 8848 10912
rect 8912 10848 8928 10912
rect 8992 10848 9008 10912
rect 9072 10848 9088 10912
rect 9152 10848 9160 10912
rect 8840 9824 9160 10848
rect 9446 10709 9506 12547
rect 9443 10708 9509 10709
rect 9443 10644 9444 10708
rect 9508 10644 9509 10708
rect 9443 10643 9509 10644
rect 9443 10436 9509 10437
rect 9443 10372 9444 10436
rect 9508 10372 9509 10436
rect 9443 10371 9509 10372
rect 8840 9760 8848 9824
rect 8912 9760 8928 9824
rect 8992 9760 9008 9824
rect 9072 9760 9088 9824
rect 9152 9760 9160 9824
rect 8840 8736 9160 9760
rect 8840 8672 8848 8736
rect 8912 8672 8928 8736
rect 8992 8672 9008 8736
rect 9072 8672 9088 8736
rect 9152 8672 9160 8736
rect 8840 7648 9160 8672
rect 9446 7717 9506 10371
rect 9630 9757 9690 14315
rect 9814 12205 9874 14995
rect 9811 12204 9877 12205
rect 9811 12140 9812 12204
rect 9876 12140 9877 12204
rect 9811 12139 9877 12140
rect 9811 12068 9877 12069
rect 9811 12004 9812 12068
rect 9876 12004 9877 12068
rect 9811 12003 9877 12004
rect 9627 9756 9693 9757
rect 9627 9692 9628 9756
rect 9692 9692 9693 9756
rect 9627 9691 9693 9692
rect 9627 8260 9693 8261
rect 9627 8196 9628 8260
rect 9692 8196 9693 8260
rect 9627 8195 9693 8196
rect 9630 7989 9690 8195
rect 9814 8125 9874 12003
rect 9998 10709 10058 16355
rect 10179 15060 10245 15061
rect 10179 14996 10180 15060
rect 10244 14996 10245 15060
rect 10179 14995 10245 14996
rect 10182 10981 10242 14995
rect 10363 14244 10429 14245
rect 10363 14180 10364 14244
rect 10428 14180 10429 14244
rect 10363 14179 10429 14180
rect 10366 12341 10426 14179
rect 10363 12340 10429 12341
rect 10363 12276 10364 12340
rect 10428 12276 10429 12340
rect 10363 12275 10429 12276
rect 10366 12069 10426 12275
rect 10363 12068 10429 12069
rect 10363 12004 10364 12068
rect 10428 12004 10429 12068
rect 10363 12003 10429 12004
rect 10550 11522 10610 17307
rect 10366 11462 10610 11522
rect 10814 16896 11134 17920
rect 10814 16832 10822 16896
rect 10886 16832 10902 16896
rect 10966 16832 10982 16896
rect 11046 16832 11062 16896
rect 11126 16832 11134 16896
rect 10814 15808 11134 16832
rect 10814 15744 10822 15808
rect 10886 15744 10902 15808
rect 10966 15744 10982 15808
rect 11046 15744 11062 15808
rect 11126 15744 11134 15808
rect 10814 14720 11134 15744
rect 11283 15196 11349 15197
rect 11283 15132 11284 15196
rect 11348 15132 11349 15196
rect 11283 15131 11349 15132
rect 10814 14656 10822 14720
rect 10886 14656 10902 14720
rect 10966 14656 10982 14720
rect 11046 14656 11062 14720
rect 11126 14656 11134 14720
rect 10814 13632 11134 14656
rect 11286 14245 11346 15131
rect 11283 14244 11349 14245
rect 11283 14180 11284 14244
rect 11348 14180 11349 14244
rect 11283 14179 11349 14180
rect 11283 13700 11349 13701
rect 11283 13636 11284 13700
rect 11348 13636 11349 13700
rect 11283 13635 11349 13636
rect 10814 13568 10822 13632
rect 10886 13568 10902 13632
rect 10966 13568 10982 13632
rect 11046 13568 11062 13632
rect 11126 13568 11134 13632
rect 10814 12544 11134 13568
rect 10814 12480 10822 12544
rect 10886 12480 10902 12544
rect 10966 12480 10982 12544
rect 11046 12480 11062 12544
rect 11126 12480 11134 12544
rect 10179 10980 10245 10981
rect 10179 10916 10180 10980
rect 10244 10916 10245 10980
rect 10179 10915 10245 10916
rect 10366 10842 10426 11462
rect 10182 10782 10426 10842
rect 10814 11456 11134 12480
rect 10814 11392 10822 11456
rect 10886 11392 10902 11456
rect 10966 11392 10982 11456
rect 11046 11392 11062 11456
rect 11126 11392 11134 11456
rect 9995 10708 10061 10709
rect 9995 10644 9996 10708
rect 10060 10644 10061 10708
rect 9995 10643 10061 10644
rect 10182 10437 10242 10782
rect 10363 10708 10429 10709
rect 10363 10644 10364 10708
rect 10428 10644 10429 10708
rect 10363 10643 10429 10644
rect 10179 10436 10245 10437
rect 10179 10372 10180 10436
rect 10244 10372 10245 10436
rect 10179 10371 10245 10372
rect 9995 10028 10061 10029
rect 9995 9964 9996 10028
rect 10060 9964 10061 10028
rect 9995 9963 10061 9964
rect 9811 8124 9877 8125
rect 9811 8060 9812 8124
rect 9876 8060 9877 8124
rect 9811 8059 9877 8060
rect 9627 7988 9693 7989
rect 9627 7924 9628 7988
rect 9692 7924 9693 7988
rect 9627 7923 9693 7924
rect 9627 7852 9693 7853
rect 9627 7788 9628 7852
rect 9692 7788 9693 7852
rect 9627 7787 9693 7788
rect 9443 7716 9509 7717
rect 9443 7652 9444 7716
rect 9508 7652 9509 7716
rect 9443 7651 9509 7652
rect 8840 7584 8848 7648
rect 8912 7584 8928 7648
rect 8992 7584 9008 7648
rect 9072 7584 9088 7648
rect 9152 7584 9160 7648
rect 8840 6560 9160 7584
rect 9259 7036 9325 7037
rect 9259 6972 9260 7036
rect 9324 6972 9325 7036
rect 9259 6971 9325 6972
rect 8840 6496 8848 6560
rect 8912 6496 8928 6560
rect 8992 6496 9008 6560
rect 9072 6496 9088 6560
rect 9152 6496 9160 6560
rect 8840 5472 9160 6496
rect 8840 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9008 5472
rect 9072 5408 9088 5472
rect 9152 5408 9160 5472
rect 8707 4860 8773 4861
rect 8707 4796 8708 4860
rect 8772 4796 8773 4860
rect 8707 4795 8773 4796
rect 8840 4384 9160 5408
rect 9262 5405 9322 6971
rect 9630 6930 9690 7787
rect 9998 7445 10058 9963
rect 10179 9756 10245 9757
rect 10179 9692 10180 9756
rect 10244 9692 10245 9756
rect 10179 9691 10245 9692
rect 9995 7444 10061 7445
rect 9995 7380 9996 7444
rect 10060 7380 10061 7444
rect 9995 7379 10061 7380
rect 9811 7172 9877 7173
rect 9811 7108 9812 7172
rect 9876 7108 9877 7172
rect 9811 7107 9877 7108
rect 9446 6870 9690 6930
rect 9259 5404 9325 5405
rect 9259 5340 9260 5404
rect 9324 5340 9325 5404
rect 9259 5339 9325 5340
rect 8840 4320 8848 4384
rect 8912 4320 8928 4384
rect 8992 4320 9008 4384
rect 9072 4320 9088 4384
rect 9152 4320 9160 4384
rect 8707 4316 8773 4317
rect 8707 4252 8708 4316
rect 8772 4252 8773 4316
rect 8707 4251 8773 4252
rect 8710 3773 8770 4251
rect 8707 3772 8773 3773
rect 8707 3708 8708 3772
rect 8772 3708 8773 3772
rect 8707 3707 8773 3708
rect 8523 3364 8589 3365
rect 8523 3300 8524 3364
rect 8588 3300 8589 3364
rect 8523 3299 8589 3300
rect 8840 3296 9160 4320
rect 8840 3232 8848 3296
rect 8912 3232 8928 3296
rect 8992 3232 9008 3296
rect 9072 3232 9088 3296
rect 9152 3232 9160 3296
rect 7787 2276 7853 2277
rect 7787 2212 7788 2276
rect 7852 2212 7853 2276
rect 7787 2211 7853 2212
rect 8155 2276 8221 2277
rect 8155 2212 8156 2276
rect 8220 2212 8221 2276
rect 8155 2211 8221 2212
rect 6866 1600 6874 1664
rect 6938 1600 6954 1664
rect 7018 1600 7034 1664
rect 7098 1600 7114 1664
rect 7178 1600 7186 1664
rect 6866 1040 7186 1600
rect 8158 1461 8218 2211
rect 8840 2208 9160 3232
rect 9262 3229 9322 5339
rect 9259 3228 9325 3229
rect 9259 3164 9260 3228
rect 9324 3164 9325 3228
rect 9259 3163 9325 3164
rect 8840 2144 8848 2208
rect 8912 2144 8928 2208
rect 8992 2144 9008 2208
rect 9072 2144 9088 2208
rect 9152 2144 9160 2208
rect 8155 1460 8221 1461
rect 8155 1396 8156 1460
rect 8220 1396 8221 1460
rect 8155 1395 8221 1396
rect 8840 1120 9160 2144
rect 9446 2141 9506 6870
rect 9627 5948 9693 5949
rect 9627 5884 9628 5948
rect 9692 5884 9693 5948
rect 9627 5883 9693 5884
rect 9630 5541 9690 5883
rect 9627 5540 9693 5541
rect 9627 5476 9628 5540
rect 9692 5476 9693 5540
rect 9627 5475 9693 5476
rect 9630 4725 9690 5475
rect 9814 4861 9874 7107
rect 10182 6930 10242 9691
rect 9998 6870 10242 6930
rect 9811 4860 9877 4861
rect 9811 4796 9812 4860
rect 9876 4796 9877 4860
rect 9811 4795 9877 4796
rect 9627 4724 9693 4725
rect 9627 4660 9628 4724
rect 9692 4660 9693 4724
rect 9627 4659 9693 4660
rect 9811 4724 9877 4725
rect 9811 4660 9812 4724
rect 9876 4660 9877 4724
rect 9811 4659 9877 4660
rect 9814 2549 9874 4659
rect 9998 3909 10058 6870
rect 10179 6764 10245 6765
rect 10179 6700 10180 6764
rect 10244 6700 10245 6764
rect 10179 6699 10245 6700
rect 9995 3908 10061 3909
rect 9995 3844 9996 3908
rect 10060 3844 10061 3908
rect 9995 3843 10061 3844
rect 10182 2685 10242 6699
rect 10366 5541 10426 10643
rect 10814 10368 11134 11392
rect 10814 10304 10822 10368
rect 10886 10304 10902 10368
rect 10966 10304 10982 10368
rect 11046 10304 11062 10368
rect 11126 10304 11134 10368
rect 10547 9484 10613 9485
rect 10547 9420 10548 9484
rect 10612 9420 10613 9484
rect 10547 9419 10613 9420
rect 10550 8805 10610 9419
rect 10814 9280 11134 10304
rect 11286 9621 11346 13635
rect 11470 12477 11530 18395
rect 12571 18188 12637 18189
rect 12571 18124 12572 18188
rect 12636 18124 12637 18188
rect 12571 18123 12637 18124
rect 11651 17508 11717 17509
rect 11651 17444 11652 17508
rect 11716 17444 11717 17508
rect 11651 17443 11717 17444
rect 11654 13157 11714 17443
rect 12019 16420 12085 16421
rect 12019 16356 12020 16420
rect 12084 16356 12085 16420
rect 12019 16355 12085 16356
rect 11835 16012 11901 16013
rect 11835 15948 11836 16012
rect 11900 15948 11901 16012
rect 11835 15947 11901 15948
rect 11651 13156 11717 13157
rect 11651 13092 11652 13156
rect 11716 13092 11717 13156
rect 11651 13091 11717 13092
rect 11651 13020 11717 13021
rect 11651 12956 11652 13020
rect 11716 12956 11717 13020
rect 11651 12955 11717 12956
rect 11467 12476 11533 12477
rect 11467 12412 11468 12476
rect 11532 12412 11533 12476
rect 11467 12411 11533 12412
rect 11467 12340 11533 12341
rect 11467 12276 11468 12340
rect 11532 12276 11533 12340
rect 11467 12275 11533 12276
rect 11470 11117 11530 12275
rect 11467 11116 11533 11117
rect 11467 11052 11468 11116
rect 11532 11052 11533 11116
rect 11467 11051 11533 11052
rect 11467 10980 11533 10981
rect 11467 10916 11468 10980
rect 11532 10916 11533 10980
rect 11467 10915 11533 10916
rect 11470 10706 11530 10915
rect 11654 10842 11714 12955
rect 11838 11525 11898 15947
rect 11835 11524 11901 11525
rect 11835 11460 11836 11524
rect 11900 11460 11901 11524
rect 11835 11459 11901 11460
rect 11835 10844 11901 10845
rect 11835 10842 11836 10844
rect 11654 10782 11836 10842
rect 11835 10780 11836 10782
rect 11900 10780 11901 10844
rect 11835 10779 11901 10780
rect 11470 10646 11714 10706
rect 11467 10436 11533 10437
rect 11467 10372 11468 10436
rect 11532 10372 11533 10436
rect 11467 10371 11533 10372
rect 11283 9620 11349 9621
rect 11283 9556 11284 9620
rect 11348 9556 11349 9620
rect 11283 9555 11349 9556
rect 11470 9482 11530 10371
rect 11654 9621 11714 10646
rect 11838 10434 11898 10779
rect 12022 10573 12082 16355
rect 12387 15196 12453 15197
rect 12387 15132 12388 15196
rect 12452 15132 12453 15196
rect 12387 15131 12453 15132
rect 12203 14652 12269 14653
rect 12203 14588 12204 14652
rect 12268 14588 12269 14652
rect 12203 14587 12269 14588
rect 12019 10572 12085 10573
rect 12019 10508 12020 10572
rect 12084 10508 12085 10572
rect 12019 10507 12085 10508
rect 11838 10374 12082 10434
rect 11651 9620 11717 9621
rect 11651 9556 11652 9620
rect 11716 9556 11717 9620
rect 11651 9555 11717 9556
rect 10814 9216 10822 9280
rect 10886 9216 10902 9280
rect 10966 9216 10982 9280
rect 11046 9216 11062 9280
rect 11126 9216 11134 9280
rect 10547 8804 10613 8805
rect 10547 8740 10548 8804
rect 10612 8740 10613 8804
rect 10547 8739 10613 8740
rect 10363 5540 10429 5541
rect 10363 5476 10364 5540
rect 10428 5476 10429 5540
rect 10363 5475 10429 5476
rect 10363 4996 10429 4997
rect 10363 4932 10364 4996
rect 10428 4932 10429 4996
rect 10363 4931 10429 4932
rect 10179 2684 10245 2685
rect 10179 2620 10180 2684
rect 10244 2620 10245 2684
rect 10179 2619 10245 2620
rect 9811 2548 9877 2549
rect 9811 2484 9812 2548
rect 9876 2484 9877 2548
rect 9811 2483 9877 2484
rect 10366 2141 10426 4931
rect 10550 3093 10610 8739
rect 10814 8192 11134 9216
rect 10814 8128 10822 8192
rect 10886 8128 10902 8192
rect 10966 8128 10982 8192
rect 11046 8128 11062 8192
rect 11126 8128 11134 8192
rect 10814 7104 11134 8128
rect 11286 9422 11530 9482
rect 11286 7173 11346 9422
rect 11651 8396 11717 8397
rect 11651 8332 11652 8396
rect 11716 8332 11717 8396
rect 11651 8331 11717 8332
rect 11467 7852 11533 7853
rect 11467 7788 11468 7852
rect 11532 7788 11533 7852
rect 11467 7787 11533 7788
rect 11283 7172 11349 7173
rect 11283 7108 11284 7172
rect 11348 7108 11349 7172
rect 11283 7107 11349 7108
rect 10814 7040 10822 7104
rect 10886 7040 10902 7104
rect 10966 7040 10982 7104
rect 11046 7040 11062 7104
rect 11126 7040 11134 7104
rect 10814 6016 11134 7040
rect 11283 6900 11349 6901
rect 11283 6836 11284 6900
rect 11348 6836 11349 6900
rect 11283 6835 11349 6836
rect 10814 5952 10822 6016
rect 10886 5952 10902 6016
rect 10966 5952 10982 6016
rect 11046 5952 11062 6016
rect 11126 5952 11134 6016
rect 10814 4928 11134 5952
rect 10814 4864 10822 4928
rect 10886 4864 10902 4928
rect 10966 4864 10982 4928
rect 11046 4864 11062 4928
rect 11126 4864 11134 4928
rect 10814 3840 11134 4864
rect 11286 4725 11346 6835
rect 11470 6085 11530 7787
rect 11467 6084 11533 6085
rect 11467 6020 11468 6084
rect 11532 6020 11533 6084
rect 11467 6019 11533 6020
rect 11467 5540 11533 5541
rect 11467 5476 11468 5540
rect 11532 5476 11533 5540
rect 11467 5475 11533 5476
rect 11283 4724 11349 4725
rect 11283 4660 11284 4724
rect 11348 4660 11349 4724
rect 11283 4659 11349 4660
rect 10814 3776 10822 3840
rect 10886 3776 10902 3840
rect 10966 3776 10982 3840
rect 11046 3776 11062 3840
rect 11126 3776 11134 3840
rect 10547 3092 10613 3093
rect 10547 3028 10548 3092
rect 10612 3028 10613 3092
rect 10547 3027 10613 3028
rect 10814 2752 11134 3776
rect 10814 2688 10822 2752
rect 10886 2688 10902 2752
rect 10966 2688 10982 2752
rect 11046 2688 11062 2752
rect 11126 2688 11134 2752
rect 9443 2140 9509 2141
rect 9443 2076 9444 2140
rect 9508 2076 9509 2140
rect 9443 2075 9509 2076
rect 10363 2140 10429 2141
rect 10363 2076 10364 2140
rect 10428 2076 10429 2140
rect 10363 2075 10429 2076
rect 8840 1056 8848 1120
rect 8912 1056 8928 1120
rect 8992 1056 9008 1120
rect 9072 1056 9088 1120
rect 9152 1056 9160 1120
rect 8840 1040 9160 1056
rect 9446 645 9506 2075
rect 10814 1664 11134 2688
rect 11470 1733 11530 5475
rect 11654 3773 11714 8331
rect 11835 8124 11901 8125
rect 11835 8060 11836 8124
rect 11900 8060 11901 8124
rect 11835 8059 11901 8060
rect 11838 4861 11898 8059
rect 12022 4997 12082 10374
rect 12206 8397 12266 14587
rect 12390 12069 12450 15131
rect 12387 12068 12453 12069
rect 12387 12004 12388 12068
rect 12452 12004 12453 12068
rect 12387 12003 12453 12004
rect 12387 11932 12453 11933
rect 12387 11868 12388 11932
rect 12452 11868 12453 11932
rect 12387 11867 12453 11868
rect 12203 8396 12269 8397
rect 12203 8332 12204 8396
rect 12268 8332 12269 8396
rect 12203 8331 12269 8332
rect 12390 8125 12450 11867
rect 12574 8669 12634 18123
rect 12788 17440 13108 18464
rect 12788 17376 12796 17440
rect 12860 17376 12876 17440
rect 12940 17376 12956 17440
rect 13020 17376 13036 17440
rect 13100 17376 13108 17440
rect 12788 16352 13108 17376
rect 14762 22336 15082 22896
rect 16619 22540 16685 22541
rect 16619 22476 16620 22540
rect 16684 22476 16685 22540
rect 16619 22475 16685 22476
rect 14762 22272 14770 22336
rect 14834 22272 14850 22336
rect 14914 22272 14930 22336
rect 14994 22272 15010 22336
rect 15074 22272 15082 22336
rect 14762 21248 15082 22272
rect 14762 21184 14770 21248
rect 14834 21184 14850 21248
rect 14914 21184 14930 21248
rect 14994 21184 15010 21248
rect 15074 21184 15082 21248
rect 14762 20160 15082 21184
rect 14762 20096 14770 20160
rect 14834 20096 14850 20160
rect 14914 20096 14930 20160
rect 14994 20096 15010 20160
rect 15074 20096 15082 20160
rect 14762 19072 15082 20096
rect 14762 19008 14770 19072
rect 14834 19008 14850 19072
rect 14914 19008 14930 19072
rect 14994 19008 15010 19072
rect 15074 19008 15082 19072
rect 14762 17984 15082 19008
rect 14762 17920 14770 17984
rect 14834 17920 14850 17984
rect 14914 17920 14930 17984
rect 14994 17920 15010 17984
rect 15074 17920 15082 17984
rect 14043 17100 14109 17101
rect 14043 17036 14044 17100
rect 14108 17036 14109 17100
rect 14043 17035 14109 17036
rect 12788 16288 12796 16352
rect 12860 16288 12876 16352
rect 12940 16288 12956 16352
rect 13020 16288 13036 16352
rect 13100 16288 13108 16352
rect 12788 15264 13108 16288
rect 13859 15468 13925 15469
rect 13859 15404 13860 15468
rect 13924 15404 13925 15468
rect 13859 15403 13925 15404
rect 12788 15200 12796 15264
rect 12860 15200 12876 15264
rect 12940 15200 12956 15264
rect 13020 15200 13036 15264
rect 13100 15200 13108 15264
rect 12788 14176 13108 15200
rect 13675 14788 13741 14789
rect 13675 14724 13676 14788
rect 13740 14724 13741 14788
rect 13675 14723 13741 14724
rect 13491 14516 13557 14517
rect 13491 14452 13492 14516
rect 13556 14452 13557 14516
rect 13491 14451 13557 14452
rect 13307 14244 13373 14245
rect 13307 14180 13308 14244
rect 13372 14180 13373 14244
rect 13307 14179 13373 14180
rect 12788 14112 12796 14176
rect 12860 14112 12876 14176
rect 12940 14112 12956 14176
rect 13020 14112 13036 14176
rect 13100 14112 13108 14176
rect 12788 13088 13108 14112
rect 13169 13564 13235 13565
rect 13169 13500 13170 13564
rect 13234 13500 13235 13564
rect 13169 13499 13235 13500
rect 12788 13024 12796 13088
rect 12860 13024 12876 13088
rect 12940 13024 12956 13088
rect 13020 13024 13036 13088
rect 13100 13024 13108 13088
rect 12788 12000 13108 13024
rect 12788 11936 12796 12000
rect 12860 11936 12876 12000
rect 12940 11936 12956 12000
rect 13020 11936 13036 12000
rect 13100 11936 13108 12000
rect 12788 10912 13108 11936
rect 13172 11525 13232 13499
rect 13169 11524 13235 11525
rect 13169 11460 13170 11524
rect 13234 11460 13235 11524
rect 13169 11459 13235 11460
rect 12788 10848 12796 10912
rect 12860 10848 12876 10912
rect 12940 10848 12956 10912
rect 13020 10848 13036 10912
rect 13100 10848 13108 10912
rect 12788 9824 13108 10848
rect 12788 9760 12796 9824
rect 12860 9760 12876 9824
rect 12940 9760 12956 9824
rect 13020 9760 13036 9824
rect 13100 9760 13108 9824
rect 12788 8736 13108 9760
rect 13310 9485 13370 14179
rect 13307 9484 13373 9485
rect 13307 9420 13308 9484
rect 13372 9420 13373 9484
rect 13307 9419 13373 9420
rect 12788 8672 12796 8736
rect 12860 8672 12876 8736
rect 12940 8672 12956 8736
rect 13020 8672 13036 8736
rect 13100 8672 13108 8736
rect 12571 8668 12637 8669
rect 12571 8604 12572 8668
rect 12636 8604 12637 8668
rect 12571 8603 12637 8604
rect 12387 8124 12453 8125
rect 12387 8060 12388 8124
rect 12452 8060 12453 8124
rect 12387 8059 12453 8060
rect 12387 7988 12453 7989
rect 12387 7924 12388 7988
rect 12452 7924 12453 7988
rect 12387 7923 12453 7924
rect 12203 7852 12269 7853
rect 12203 7788 12204 7852
rect 12268 7788 12269 7852
rect 12203 7787 12269 7788
rect 12206 5541 12266 7787
rect 12390 6357 12450 7923
rect 12571 7852 12637 7853
rect 12571 7788 12572 7852
rect 12636 7788 12637 7852
rect 12571 7787 12637 7788
rect 12387 6356 12453 6357
rect 12387 6292 12388 6356
rect 12452 6292 12453 6356
rect 12387 6291 12453 6292
rect 12203 5540 12269 5541
rect 12203 5476 12204 5540
rect 12268 5476 12269 5540
rect 12203 5475 12269 5476
rect 12019 4996 12085 4997
rect 12019 4932 12020 4996
rect 12084 4932 12085 4996
rect 12019 4931 12085 4932
rect 12203 4996 12269 4997
rect 12203 4932 12204 4996
rect 12268 4932 12269 4996
rect 12203 4931 12269 4932
rect 11835 4860 11901 4861
rect 11835 4796 11836 4860
rect 11900 4796 11901 4860
rect 11835 4795 11901 4796
rect 12019 4724 12085 4725
rect 12019 4660 12020 4724
rect 12084 4660 12085 4724
rect 12019 4659 12085 4660
rect 12022 3909 12082 4659
rect 12019 3908 12085 3909
rect 12019 3844 12020 3908
rect 12084 3844 12085 3908
rect 12019 3843 12085 3844
rect 11651 3772 11717 3773
rect 11651 3708 11652 3772
rect 11716 3708 11717 3772
rect 11651 3707 11717 3708
rect 12206 2685 12266 4931
rect 12390 2821 12450 6291
rect 12387 2820 12453 2821
rect 12387 2756 12388 2820
rect 12452 2756 12453 2820
rect 12387 2755 12453 2756
rect 12203 2684 12269 2685
rect 12203 2620 12204 2684
rect 12268 2620 12269 2684
rect 12203 2619 12269 2620
rect 12390 2141 12450 2755
rect 12387 2140 12453 2141
rect 12387 2076 12388 2140
rect 12452 2076 12453 2140
rect 12387 2075 12453 2076
rect 12574 1733 12634 7787
rect 12788 7648 13108 8672
rect 13307 8668 13373 8669
rect 13307 8604 13308 8668
rect 13372 8604 13373 8668
rect 13307 8603 13373 8604
rect 12788 7584 12796 7648
rect 12860 7584 12876 7648
rect 12940 7584 12956 7648
rect 13020 7584 13036 7648
rect 13100 7584 13108 7648
rect 12788 6560 13108 7584
rect 12788 6496 12796 6560
rect 12860 6496 12876 6560
rect 12940 6496 12956 6560
rect 13020 6496 13036 6560
rect 13100 6496 13108 6560
rect 12788 5472 13108 6496
rect 12788 5408 12796 5472
rect 12860 5408 12876 5472
rect 12940 5408 12956 5472
rect 13020 5408 13036 5472
rect 13100 5408 13108 5472
rect 12788 4384 13108 5408
rect 13310 4725 13370 8603
rect 13494 4861 13554 14451
rect 13678 6493 13738 14723
rect 13862 11797 13922 15403
rect 14046 12885 14106 17035
rect 14762 16896 15082 17920
rect 14762 16832 14770 16896
rect 14834 16832 14850 16896
rect 14914 16832 14930 16896
rect 14994 16832 15010 16896
rect 15074 16832 15082 16896
rect 14762 15808 15082 16832
rect 14762 15744 14770 15808
rect 14834 15744 14850 15808
rect 14914 15744 14930 15808
rect 14994 15744 15010 15808
rect 15074 15744 15082 15808
rect 14762 14720 15082 15744
rect 15883 15604 15949 15605
rect 15883 15540 15884 15604
rect 15948 15540 15949 15604
rect 15883 15539 15949 15540
rect 15515 15060 15581 15061
rect 15515 14996 15516 15060
rect 15580 14996 15581 15060
rect 15515 14995 15581 14996
rect 14762 14656 14770 14720
rect 14834 14656 14850 14720
rect 14914 14656 14930 14720
rect 14994 14656 15010 14720
rect 15074 14656 15082 14720
rect 14411 13972 14477 13973
rect 14411 13908 14412 13972
rect 14476 13908 14477 13972
rect 14411 13907 14477 13908
rect 14227 13564 14293 13565
rect 14227 13500 14228 13564
rect 14292 13500 14293 13564
rect 14227 13499 14293 13500
rect 14043 12884 14109 12885
rect 14043 12820 14044 12884
rect 14108 12820 14109 12884
rect 14043 12819 14109 12820
rect 14043 12204 14109 12205
rect 14043 12140 14044 12204
rect 14108 12140 14109 12204
rect 14043 12139 14109 12140
rect 14046 12069 14106 12139
rect 14043 12068 14109 12069
rect 14043 12004 14044 12068
rect 14108 12004 14109 12068
rect 14043 12003 14109 12004
rect 13859 11796 13925 11797
rect 13859 11732 13860 11796
rect 13924 11732 13925 11796
rect 13859 11731 13925 11732
rect 13859 11660 13925 11661
rect 13859 11596 13860 11660
rect 13924 11596 13925 11660
rect 13859 11595 13925 11596
rect 13862 8941 13922 11595
rect 14043 11524 14109 11525
rect 14043 11460 14044 11524
rect 14108 11460 14109 11524
rect 14043 11459 14109 11460
rect 14046 10845 14106 11459
rect 14043 10844 14109 10845
rect 14043 10780 14044 10844
rect 14108 10780 14109 10844
rect 14043 10779 14109 10780
rect 14230 10434 14290 13499
rect 14414 11117 14474 13907
rect 14595 13700 14661 13701
rect 14595 13636 14596 13700
rect 14660 13636 14661 13700
rect 14595 13635 14661 13636
rect 14411 11116 14477 11117
rect 14411 11052 14412 11116
rect 14476 11052 14477 11116
rect 14411 11051 14477 11052
rect 14598 10437 14658 13635
rect 14762 13632 15082 14656
rect 14762 13568 14770 13632
rect 14834 13568 14850 13632
rect 14914 13568 14930 13632
rect 14994 13568 15010 13632
rect 15074 13568 15082 13632
rect 14762 12544 15082 13568
rect 15331 13564 15397 13565
rect 15331 13500 15332 13564
rect 15396 13500 15397 13564
rect 15331 13499 15397 13500
rect 15147 13292 15213 13293
rect 15147 13228 15148 13292
rect 15212 13228 15213 13292
rect 15147 13227 15213 13228
rect 14762 12480 14770 12544
rect 14834 12480 14850 12544
rect 14914 12480 14930 12544
rect 14994 12480 15010 12544
rect 15074 12480 15082 12544
rect 14762 11456 15082 12480
rect 15150 12205 15210 13227
rect 15147 12204 15213 12205
rect 15147 12140 15148 12204
rect 15212 12140 15213 12204
rect 15147 12139 15213 12140
rect 15147 11796 15213 11797
rect 15147 11732 15148 11796
rect 15212 11732 15213 11796
rect 15147 11731 15213 11732
rect 14762 11392 14770 11456
rect 14834 11392 14850 11456
rect 14914 11392 14930 11456
rect 14994 11392 15010 11456
rect 15074 11392 15082 11456
rect 14595 10436 14661 10437
rect 14230 10374 14474 10434
rect 14043 9076 14109 9077
rect 14043 9012 14044 9076
rect 14108 9012 14109 9076
rect 14043 9011 14109 9012
rect 13859 8940 13925 8941
rect 13859 8876 13860 8940
rect 13924 8876 13925 8940
rect 13859 8875 13925 8876
rect 13862 7853 13922 8875
rect 13859 7852 13925 7853
rect 13859 7788 13860 7852
rect 13924 7788 13925 7852
rect 13859 7787 13925 7788
rect 13675 6492 13741 6493
rect 13675 6428 13676 6492
rect 13740 6428 13741 6492
rect 13675 6427 13741 6428
rect 13859 6356 13925 6357
rect 13859 6292 13860 6356
rect 13924 6292 13925 6356
rect 13859 6291 13925 6292
rect 13675 5812 13741 5813
rect 13675 5748 13676 5812
rect 13740 5748 13741 5812
rect 13675 5747 13741 5748
rect 13491 4860 13557 4861
rect 13491 4796 13492 4860
rect 13556 4796 13557 4860
rect 13491 4795 13557 4796
rect 13307 4724 13373 4725
rect 13307 4660 13308 4724
rect 13372 4660 13373 4724
rect 13307 4659 13373 4660
rect 12788 4320 12796 4384
rect 12860 4320 12876 4384
rect 12940 4320 12956 4384
rect 13020 4320 13036 4384
rect 13100 4320 13108 4384
rect 12788 3296 13108 4320
rect 12788 3232 12796 3296
rect 12860 3232 12876 3296
rect 12940 3232 12956 3296
rect 13020 3232 13036 3296
rect 13100 3232 13108 3296
rect 12788 2208 13108 3232
rect 13494 3093 13554 4795
rect 13491 3092 13557 3093
rect 13491 3028 13492 3092
rect 13556 3028 13557 3092
rect 13491 3027 13557 3028
rect 12788 2144 12796 2208
rect 12860 2144 12876 2208
rect 12940 2144 12956 2208
rect 13020 2144 13036 2208
rect 13100 2144 13108 2208
rect 11467 1732 11533 1733
rect 11467 1668 11468 1732
rect 11532 1668 11533 1732
rect 11467 1667 11533 1668
rect 12571 1732 12637 1733
rect 12571 1668 12572 1732
rect 12636 1668 12637 1732
rect 12571 1667 12637 1668
rect 10814 1600 10822 1664
rect 10886 1600 10902 1664
rect 10966 1600 10982 1664
rect 11046 1600 11062 1664
rect 11126 1600 11134 1664
rect 10814 1040 11134 1600
rect 12788 1120 13108 2144
rect 13494 1597 13554 3027
rect 13678 1869 13738 5747
rect 13675 1868 13741 1869
rect 13675 1804 13676 1868
rect 13740 1804 13741 1868
rect 13675 1803 13741 1804
rect 13491 1596 13557 1597
rect 13491 1532 13492 1596
rect 13556 1532 13557 1596
rect 13491 1531 13557 1532
rect 12788 1056 12796 1120
rect 12860 1056 12876 1120
rect 12940 1056 12956 1120
rect 13020 1056 13036 1120
rect 13100 1056 13108 1120
rect 12788 1040 13108 1056
rect 13862 645 13922 6291
rect 14046 3637 14106 9011
rect 14414 8669 14474 10374
rect 14595 10372 14596 10436
rect 14660 10372 14661 10436
rect 14595 10371 14661 10372
rect 14762 10368 15082 11392
rect 14762 10304 14770 10368
rect 14834 10304 14850 10368
rect 14914 10304 14930 10368
rect 14994 10304 15010 10368
rect 15074 10304 15082 10368
rect 14762 9280 15082 10304
rect 14762 9216 14770 9280
rect 14834 9216 14850 9280
rect 14914 9216 14930 9280
rect 14994 9216 15010 9280
rect 15074 9216 15082 9280
rect 14411 8668 14477 8669
rect 14411 8604 14412 8668
rect 14476 8604 14477 8668
rect 14411 8603 14477 8604
rect 14411 8532 14477 8533
rect 14411 8468 14412 8532
rect 14476 8468 14477 8532
rect 14411 8467 14477 8468
rect 14227 8260 14293 8261
rect 14227 8196 14228 8260
rect 14292 8196 14293 8260
rect 14227 8195 14293 8196
rect 14230 4453 14290 8195
rect 14414 5949 14474 8467
rect 14762 8192 15082 9216
rect 14762 8128 14770 8192
rect 14834 8128 14850 8192
rect 14914 8128 14930 8192
rect 14994 8128 15010 8192
rect 15074 8128 15082 8192
rect 14762 7104 15082 8128
rect 14762 7040 14770 7104
rect 14834 7040 14850 7104
rect 14914 7040 14930 7104
rect 14994 7040 15010 7104
rect 15074 7040 15082 7104
rect 14762 6016 15082 7040
rect 14762 5952 14770 6016
rect 14834 5952 14850 6016
rect 14914 5952 14930 6016
rect 14994 5952 15010 6016
rect 15074 5952 15082 6016
rect 14411 5948 14477 5949
rect 14411 5884 14412 5948
rect 14476 5884 14477 5948
rect 14411 5883 14477 5884
rect 14762 4928 15082 5952
rect 15150 5133 15210 11731
rect 15334 6901 15394 13499
rect 15518 12885 15578 14995
rect 15699 13292 15765 13293
rect 15699 13228 15700 13292
rect 15764 13228 15765 13292
rect 15699 13227 15765 13228
rect 15515 12884 15581 12885
rect 15515 12820 15516 12884
rect 15580 12820 15581 12884
rect 15515 12819 15581 12820
rect 15515 12612 15581 12613
rect 15515 12548 15516 12612
rect 15580 12548 15581 12612
rect 15515 12547 15581 12548
rect 15331 6900 15397 6901
rect 15331 6836 15332 6900
rect 15396 6836 15397 6900
rect 15331 6835 15397 6836
rect 15331 6628 15397 6629
rect 15331 6564 15332 6628
rect 15396 6564 15397 6628
rect 15331 6563 15397 6564
rect 15147 5132 15213 5133
rect 15147 5068 15148 5132
rect 15212 5068 15213 5132
rect 15147 5067 15213 5068
rect 14762 4864 14770 4928
rect 14834 4864 14850 4928
rect 14914 4864 14930 4928
rect 14994 4864 15010 4928
rect 15074 4864 15082 4928
rect 14227 4452 14293 4453
rect 14227 4388 14228 4452
rect 14292 4388 14293 4452
rect 14227 4387 14293 4388
rect 14762 3840 15082 4864
rect 14762 3776 14770 3840
rect 14834 3776 14850 3840
rect 14914 3776 14930 3840
rect 14994 3776 15010 3840
rect 15074 3776 15082 3840
rect 14043 3636 14109 3637
rect 14043 3572 14044 3636
rect 14108 3572 14109 3636
rect 14043 3571 14109 3572
rect 14762 2752 15082 3776
rect 14762 2688 14770 2752
rect 14834 2688 14850 2752
rect 14914 2688 14930 2752
rect 14994 2688 15010 2752
rect 15074 2688 15082 2752
rect 14762 1664 15082 2688
rect 15334 2413 15394 6563
rect 15518 4181 15578 12547
rect 15702 11661 15762 13227
rect 15699 11660 15765 11661
rect 15699 11596 15700 11660
rect 15764 11596 15765 11660
rect 15699 11595 15765 11596
rect 15886 11117 15946 15539
rect 16435 14924 16501 14925
rect 16435 14860 16436 14924
rect 16500 14860 16501 14924
rect 16435 14859 16501 14860
rect 16067 13020 16133 13021
rect 16067 12956 16068 13020
rect 16132 12956 16133 13020
rect 16067 12955 16133 12956
rect 15883 11116 15949 11117
rect 15883 11052 15884 11116
rect 15948 11052 15949 11116
rect 15883 11051 15949 11052
rect 15699 10844 15765 10845
rect 15699 10780 15700 10844
rect 15764 10780 15765 10844
rect 15699 10779 15765 10780
rect 15702 9077 15762 10779
rect 15699 9076 15765 9077
rect 15699 9012 15700 9076
rect 15764 9012 15765 9076
rect 15699 9011 15765 9012
rect 16070 8533 16130 12955
rect 16251 12204 16317 12205
rect 16251 12140 16252 12204
rect 16316 12140 16317 12204
rect 16251 12139 16317 12140
rect 16067 8532 16133 8533
rect 16067 8468 16068 8532
rect 16132 8468 16133 8532
rect 16067 8467 16133 8468
rect 15699 8396 15765 8397
rect 15699 8332 15700 8396
rect 15764 8332 15765 8396
rect 15699 8331 15765 8332
rect 15702 6629 15762 8331
rect 15699 6628 15765 6629
rect 15699 6564 15700 6628
rect 15764 6564 15765 6628
rect 15699 6563 15765 6564
rect 15515 4180 15581 4181
rect 15515 4116 15516 4180
rect 15580 4116 15581 4180
rect 15515 4115 15581 4116
rect 16070 3093 16130 8467
rect 16254 6221 16314 12139
rect 16438 9893 16498 14859
rect 16435 9892 16501 9893
rect 16435 9828 16436 9892
rect 16500 9828 16501 9892
rect 16435 9827 16501 9828
rect 16622 7581 16682 22475
rect 16803 18324 16869 18325
rect 16803 18260 16804 18324
rect 16868 18260 16869 18324
rect 16803 18259 16869 18260
rect 16619 7580 16685 7581
rect 16619 7516 16620 7580
rect 16684 7516 16685 7580
rect 16619 7515 16685 7516
rect 16251 6220 16317 6221
rect 16251 6156 16252 6220
rect 16316 6156 16317 6220
rect 16251 6155 16317 6156
rect 16806 4181 16866 18259
rect 16803 4180 16869 4181
rect 16803 4116 16804 4180
rect 16868 4116 16869 4180
rect 16803 4115 16869 4116
rect 16067 3092 16133 3093
rect 16067 3028 16068 3092
rect 16132 3028 16133 3092
rect 16067 3027 16133 3028
rect 15331 2412 15397 2413
rect 15331 2348 15332 2412
rect 15396 2348 15397 2412
rect 15331 2347 15397 2348
rect 14762 1600 14770 1664
rect 14834 1600 14850 1664
rect 14914 1600 14930 1664
rect 14994 1600 15010 1664
rect 15074 1600 15082 1664
rect 14762 1040 15082 1600
rect 9443 644 9509 645
rect 9443 580 9444 644
rect 9508 580 9509 644
rect 9443 579 9509 580
rect 13859 644 13925 645
rect 13859 580 13860 644
rect 13924 580 13925 644
rect 13859 579 13925 580
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 0
transform -1 0 10304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 0
transform 1 0 15180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 0
transform -1 0 2760 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 0
transform -1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 0
transform -1 0 14996 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 0
transform 1 0 1840 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 0
transform 1 0 1656 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 0
transform 1 0 4508 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 0
transform 1 0 1380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7
timestamp 0
transform 1 0 1748 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14
timestamp 0
transform 1 0 2392 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 0
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 0
transform 1 0 4232 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 0
transform 1 0 5244 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 0
transform 1 0 5888 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 0
transform 1 0 6900 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 0
transform 1 0 7820 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 0
transform 1 0 8464 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 0
transform 1 0 9476 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 0
transform 1 0 10304 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 0
transform 1 0 11040 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 0
transform 1 0 11960 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127
timestamp 0
transform 1 0 12788 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 0
transform 1 0 13616 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 0
transform 1 0 14536 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154
timestamp 0
transform 1 0 15272 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 0
transform 1 0 15916 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 0
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 0
transform 1 0 1380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 0
transform 1 0 2300 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 0
transform 1 0 3312 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_28
timestamp 0
transform 1 0 3680 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_38
timestamp 0
transform 1 0 4600 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_44
timestamp 0
transform 1 0 5152 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 0
transform 1 0 5888 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_61
timestamp 0
transform 1 0 6716 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 0
transform 1 0 8556 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_91
timestamp 0
transform 1 0 9476 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_101
timestamp 0
transform 1 0 10396 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 0
transform 1 0 11040 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 0
transform 1 0 11960 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 0
transform 1 0 12788 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 0
transform 1 0 13616 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 0
transform 1 0 14444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 0
transform 1 0 15088 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 0
transform 1 0 15732 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 0
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 0
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_38
timestamp 0
transform 1 0 4600 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 0
transform 1 0 5152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_65
timestamp 0
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 0
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_91
timestamp 0
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 0
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_110
timestamp 0
transform 1 0 11224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 0
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 0
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 0
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_145
timestamp 0
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_152
timestamp 0
transform 1 0 15088 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 0
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_167
timestamp 0
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_12
timestamp 0
transform 1 0 2208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_32
timestamp 0
transform 1 0 4048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 0
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_66
timestamp 0
transform 1 0 7176 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_72
timestamp 0
transform 1 0 7728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 0
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 0
transform 1 0 11960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 0
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 0
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_143
timestamp 0
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_150
timestamp 0
transform 1 0 14904 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_157
timestamp 0
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 0
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_16
timestamp 0
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 0
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_39
timestamp 0
transform 1 0 4692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 0
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_101
timestamp 0
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 0
transform 1 0 11224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_119
timestamp 0
transform 1 0 12052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_127
timestamp 0
transform 1 0 12788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 0
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_145
timestamp 0
transform 1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_152
timestamp 0
transform 1 0 15088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_159
timestamp 0
transform 1 0 15732 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_167
timestamp 0
transform 1 0 16468 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_10
timestamp 0
transform 1 0 2024 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 0
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 0
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_61
timestamp 0
transform 1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 0
transform 1 0 9108 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 0
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_119
timestamp 0
transform 1 0 12052 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 0
transform 1 0 12788 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_134
timestamp 0
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_143
timestamp 0
transform 1 0 14260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_151
timestamp 0
transform 1 0 14996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_159
timestamp 0
transform 1 0 15732 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 0
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_10
timestamp 0
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 0
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_39
timestamp 0
transform 1 0 4692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_73
timestamp 0
transform 1 0 7820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 0
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_92
timestamp 0
transform 1 0 9568 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_100
timestamp 0
transform 1 0 10304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_130
timestamp 0
transform 1 0 13064 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 0
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 0
transform 1 0 14536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_155
timestamp 0
transform 1 0 15364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 0
transform 1 0 16100 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_167
timestamp 0
transform 1 0 16468 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_8
timestamp 0
transform 1 0 1840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_28
timestamp 0
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 0
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_66
timestamp 0
transform 1 0 7176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_94
timestamp 0
transform 1 0 9752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_119
timestamp 0
transform 1 0 12052 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_147
timestamp 0
transform 1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 0
transform 1 0 14996 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_158
timestamp 0
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 0
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 0
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 0
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_119
timestamp 0
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_123
timestamp 0
transform 1 0 12420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 0
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 0
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_146
timestamp 0
transform 1 0 14536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_155
timestamp 0
transform 1 0 15364 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_164
timestamp 0
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_25
timestamp 0
transform 1 0 3404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 0
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_64
timestamp 0
transform 1 0 6992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_84
timestamp 0
transform 1 0 8832 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 0
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 0
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 0
transform 1 0 13892 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_149
timestamp 0
transform 1 0 14812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp 0
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 0
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 0
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 0
transform 1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 0
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_89
timestamp 0
transform 1 0 9292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_129
timestamp 0
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 0
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_147
timestamp 0
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_157
timestamp 0
transform 1 0 15548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 0
transform 1 0 16192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 0
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_28
timestamp 0
transform 1 0 3680 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 0
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 0
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_121
timestamp 0
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_145
timestamp 0
transform 1 0 14444 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_151
timestamp 0
transform 1 0 14996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp 0
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 0
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 0
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_39
timestamp 0
transform 1 0 4692 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 0
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_94
timestamp 0
transform 1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_100
timestamp 0
transform 1 0 10304 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_121
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 0
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_148
timestamp 0
transform 1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_158
timestamp 0
transform 1 0 15640 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_166
timestamp 0
transform 1 0 16376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_25
timestamp 0
transform 1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_49
timestamp 0
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_77
timestamp 0
transform 1 0 8188 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_83
timestamp 0
transform 1 0 8740 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 0
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 0
transform 1 0 12972 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 0
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 0
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 0
transform 1 0 15364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 0
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 0
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 0
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_36
timestamp 0
transform 1 0 4416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_60
timestamp 0
transform 1 0 6624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 0
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_129
timestamp 0
transform 1 0 12972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 0
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 0
transform 1 0 14720 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_158
timestamp 0
transform 1 0 15640 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_166
timestamp 0
transform 1 0 16376 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_14
timestamp 0
transform 1 0 2392 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_39
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 0
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_60
timestamp 0
transform 1 0 6624 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_84
timestamp 0
transform 1 0 8832 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 0
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_129
timestamp 0
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_149
timestamp 0
transform 1 0 14812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 0
transform 1 0 15732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 0
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 0
transform 1 0 4048 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 0
transform 1 0 6256 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 0
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_125
timestamp 0
transform 1 0 12604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 0
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 0
transform 1 0 14996 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_162
timestamp 0
transform 1 0 16008 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_11
timestamp 0
transform 1 0 2116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_36
timestamp 0
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 0
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_67
timestamp 0
transform 1 0 7268 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_97
timestamp 0
transform 1 0 10028 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 0
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_129
timestamp 0
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_141
timestamp 0
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 0
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 0
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 0
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 0
transform 1 0 4048 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_56
timestamp 0
transform 1 0 6256 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 0
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_101
timestamp 0
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 0
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 0
transform 1 0 14720 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_158
timestamp 0
transform 1 0 15640 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_166
timestamp 0
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_40
timestamp 0
transform 1 0 4784 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 0
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_75
timestamp 0
transform 1 0 8004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 0
transform 1 0 10212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 0
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_129
timestamp 0
transform 1 0 12972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 0
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 0
transform 1 0 14996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 0
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 0
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_50
timestamp 0
transform 1 0 5704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_58
timestamp 0
transform 1 0 6440 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 0
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_89
timestamp 0
transform 1 0 9292 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_129
timestamp 0
transform 1 0 12972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 0
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_147
timestamp 0
transform 1 0 14628 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_157
timestamp 0
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 0
transform 1 0 16192 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_16
timestamp 0
transform 1 0 2576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp 0
transform 1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 0
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_67
timestamp 0
transform 1 0 7268 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_97
timestamp 0
transform 1 0 10028 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_101
timestamp 0
transform 1 0 10396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 0
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_122
timestamp 0
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 0
transform 1 0 13524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_145
timestamp 0
transform 1 0 14444 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 0
transform 1 0 14996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 0
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 0
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 0
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_49
timestamp 0
transform 1 0 5612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_56
timestamp 0
transform 1 0 6256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 0
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_120
timestamp 0
transform 1 0 12144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 0
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_147
timestamp 0
transform 1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 0
transform 1 0 15272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 0
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_167
timestamp 0
transform 1 0 16468 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_12
timestamp 0
transform 1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_36
timestamp 0
transform 1 0 4416 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_45
timestamp 0
transform 1 0 5244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 0
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_93
timestamp 0
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 0
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_120
timestamp 0
transform 1 0 12144 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_130
timestamp 0
transform 1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_134
timestamp 0
transform 1 0 13432 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 0
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 0
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 0
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 0
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_33
timestamp 0
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_50
timestamp 0
transform 1 0 5704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 0
transform 1 0 7544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_78
timestamp 0
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_95
timestamp 0
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_108
timestamp 0
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_118
timestamp 0
transform 1 0 11960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 0
transform 1 0 12880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 0
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 0
transform 1 0 14352 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_151
timestamp 0
transform 1 0 14996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_158
timestamp 0
transform 1 0 15640 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_166
timestamp 0
transform 1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_11
timestamp 0
transform 1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 0
transform 1 0 4048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 0
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_67
timestamp 0
transform 1 0 7268 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_95
timestamp 0
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 0
transform 1 0 10856 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_119
timestamp 0
transform 1 0 12052 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_126
timestamp 0
transform 1 0 12696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_133
timestamp 0
transform 1 0 13340 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_140
timestamp 0
transform 1 0 13984 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 0
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 0
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 0
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 0
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_34
timestamp 0
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_78
timestamp 0
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_91
timestamp 0
transform 1 0 9476 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 0
transform 1 0 10396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_111
timestamp 0
transform 1 0 11316 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_118
timestamp 0
transform 1 0 11960 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 0
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_132
timestamp 0
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_147
timestamp 0
transform 1 0 14628 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_155
timestamp 0
transform 1 0 15364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_160
timestamp 0
transform 1 0 15824 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_10
timestamp 0
transform 1 0 2024 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_32
timestamp 0
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 0
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_67
timestamp 0
transform 1 0 7268 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_73
timestamp 0
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 0
transform 1 0 9292 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 0
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 0
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_116
timestamp 0
transform 1 0 11776 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_123
timestamp 0
transform 1 0 12420 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_135
timestamp 0
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_147
timestamp 0
transform 1 0 14628 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_153
timestamp 0
transform 1 0 15180 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_157
timestamp 0
transform 1 0 15548 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 0
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 0
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 0
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_33
timestamp 0
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_41
timestamp 0
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_65
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_73
timestamp 0
transform 1 0 7820 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 0
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_109
timestamp 0
transform 1 0 11132 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_116
timestamp 0
transform 1 0 11776 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_128
timestamp 0
transform 1 0 12880 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_25
timestamp 0
transform 1 0 3404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_45
timestamp 0
transform 1 0 5244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 0
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_64
timestamp 0
transform 1 0 6992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_74
timestamp 0
transform 1 0 7912 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 0
transform 1 0 8648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_89
timestamp 0
transform 1 0 9292 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_96
timestamp 0
transform 1 0 9936 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_100
timestamp 0
transform 1 0 10304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 0
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 0
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 0
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 0
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 0
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_33
timestamp 0
transform 1 0 4140 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_50
timestamp 0
transform 1 0 5704 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_54
timestamp 0
transform 1 0 6072 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 0
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_71
timestamp 0
transform 1 0 7636 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 0
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 0
transform 1 0 9200 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_95
timestamp 0
transform 1 0 9844 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_107
timestamp 0
transform 1 0 10948 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_119
timestamp 0
transform 1 0 12052 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_131
timestamp 0
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 0
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_165
timestamp 0
transform 1 0 16284 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 0
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_24
timestamp 0
transform 1 0 3312 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_28
timestamp 0
transform 1 0 3680 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_45
timestamp 0
transform 1 0 5244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 0
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_63
timestamp 0
transform 1 0 6900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_71
timestamp 0
transform 1 0 7636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_78
timestamp 0
transform 1 0 8280 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_85
timestamp 0
transform 1 0 8924 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 0
transform 1 0 9568 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 0
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 0
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 0
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_10
timestamp 0
transform 1 0 2024 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_14
timestamp 0
transform 1 0 2392 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 0
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_37
timestamp 0
transform 1 0 4508 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_51
timestamp 0
transform 1 0 5796 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_60
timestamp 0
transform 1 0 6624 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_64
timestamp 0
transform 1 0 6992 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_68
timestamp 0
transform 1 0 7360 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_75
timestamp 0
transform 1 0 8004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 0
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 0
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 0
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 0
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 0
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_165
timestamp 0
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_11
timestamp 0
transform 1 0 2116 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_22
timestamp 0
transform 1 0 3128 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_31
timestamp 0
transform 1 0 3956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 0
transform 1 0 4692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 0
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 0
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_60
timestamp 0
transform 1 0 6624 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_67
timestamp 0
transform 1 0 7268 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_79
timestamp 0
transform 1 0 8372 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_91
timestamp 0
transform 1 0 9476 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_103
timestamp 0
transform 1 0 10580 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 0
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 0
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 0
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 0
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 0
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_8
timestamp 0
transform 1 0 1840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_15
timestamp 0
transform 1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_19
timestamp 0
transform 1 0 2852 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 0
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_33
timestamp 0
transform 1 0 4140 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_40
timestamp 0
transform 1 0 4784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 0
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_54
timestamp 0
transform 1 0 6072 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_61
timestamp 0
transform 1 0 6716 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_73
timestamp 0
transform 1 0 7820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_81
timestamp 0
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 0
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 0
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 0
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 0
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 0
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_165
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_6
timestamp 0
transform 1 0 1656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 0
transform 1 0 2392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_22
timestamp 0
transform 1 0 3128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_30
timestamp 0
transform 1 0 3864 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_35
timestamp 0
transform 1 0 4324 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_39
timestamp 0
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_44
timestamp 0
transform 1 0 5152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 0
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 0
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 0
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 0
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 0
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 0
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 0
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 0
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 0
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 0
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 0
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 0
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_3
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_8
timestamp 0
transform 1 0 1840 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_16
timestamp 0
transform 1 0 2576 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 0
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_32
timestamp 0
transform 1 0 4048 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_39
timestamp 0
transform 1 0 4692 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_51
timestamp 0
transform 1 0 5796 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_63
timestamp 0
transform 1 0 6900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_75
timestamp 0
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 0
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 0
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 0
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 0
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 0
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 0
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_165
timestamp 0
transform 1 0 16284 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_8
timestamp 0
transform 1 0 1840 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_16
timestamp 0
transform 1 0 2576 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_23
timestamp 0
transform 1 0 3220 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_30
timestamp 0
transform 1 0 3864 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_42
timestamp 0
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 0
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 0
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 0
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 0
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 0
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 0
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 0
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 0
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 0
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 0
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 0
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_7
timestamp 0
transform 1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_14
timestamp 0
transform 1 0 2392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 0
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 0
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 0
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 0
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 0
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 0
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 0
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 0
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 0
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 0
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 0
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 0
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 0
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_165
timestamp 0
transform 1 0 16284 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_6
timestamp 0
transform 1 0 1656 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_10
timestamp 0
transform 1 0 2024 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_22
timestamp 0
transform 1 0 3128 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_29
timestamp 0
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_41
timestamp 0
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 0
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 0
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_81
timestamp 0
transform 1 0 8556 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_85
timestamp 0
transform 1 0 8924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_97
timestamp 0
transform 1 0 10028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 0
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 0
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_137
timestamp 0
transform 1 0 13708 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_141
timestamp 0
transform 1 0 14076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_153
timestamp 0
transform 1 0 15180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 0
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 16836 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 16836 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 0
transform -1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 0
transform -1 0 16836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 0
transform -1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 0
transform -1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 0
transform -1 0 16836 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 0
transform -1 0 16836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 0
transform -1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 0
transform -1 0 16836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 0
transform -1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 0
transform -1 0 16836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 0
transform -1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 0
transform -1 0 16836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 0
transform -1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 0
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 0
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 0
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 0
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 0
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 0
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 0
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 0
transform 1 0 3680 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 0
transform 1 0 8832 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 0
transform 1 0 13984 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _223_
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _224_
timestamp 0
transform 1 0 10672 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _225_
timestamp 0
transform 1 0 4600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _226_
timestamp 0
transform 1 0 15548 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _227_
timestamp 0
transform 1 0 13156 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 0
transform 1 0 15456 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _229_
timestamp 0
transform 1 0 14628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 0
transform 1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 0
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _232_
timestamp 0
transform 1 0 10764 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _233_
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _234_
timestamp 0
transform 1 0 8924 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _235_
timestamp 0
transform 1 0 9844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 0
transform 1 0 6992 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _237_
timestamp 0
transform 1 0 1656 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _238_
timestamp 0
transform 1 0 9844 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 0
transform 1 0 10120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _241_
timestamp 0
transform 1 0 3772 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _242_
timestamp 0
transform 1 0 2668 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _243_
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _244_
timestamp 0
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _245_
timestamp 0
transform 1 0 8924 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 0
transform 1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _247_
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _248_
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkinv_2  _249_
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _250_
timestamp 0
transform 1 0 1656 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _251_
timestamp 0
transform 1 0 12972 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _252_
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _253_
timestamp 0
transform 1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _254_
timestamp 0
transform 1 0 12512 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _255_
timestamp 0
transform 1 0 7268 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _256_
timestamp 0
transform 1 0 7912 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _257_
timestamp 0
transform 1 0 8280 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _258_
timestamp 0
transform 1 0 4876 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _259_
timestamp 0
transform 1 0 3956 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _260_
timestamp 0
transform 1 0 3496 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _261_
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _262_
timestamp 0
transform 1 0 1564 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _263_
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _264_
timestamp 0
transform 1 0 15916 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _265_
timestamp 0
transform 1 0 5612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _266_
timestamp 0
transform 1 0 5152 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _267_
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _268_
timestamp 0
transform 1 0 12420 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _269_
timestamp 0
transform 1 0 1656 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _270_
timestamp 0
transform 1 0 6164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _271_
timestamp 0
transform 1 0 14904 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _272_
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _273_
timestamp 0
transform 1 0 12328 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _274_
timestamp 0
transform 1 0 13064 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _275_
timestamp 0
transform 1 0 14352 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _276_
timestamp 0
transform 1 0 6348 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _277_
timestamp 0
transform 1 0 5612 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _278_
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _279_
timestamp 0
transform 1 0 10028 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _280_
timestamp 0
transform 1 0 4968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _281_
timestamp 0
transform 1 0 12696 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 0
transform 1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _283_
timestamp 0
transform 1 0 15548 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 0
transform 1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _285_
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _286_
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _287_
timestamp 0
transform 1 0 10028 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _288_
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp 0
transform 1 0 4048 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _290_
timestamp 0
transform 1 0 3956 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _291_
timestamp 0
transform 1 0 2852 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _293_
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _294_
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp 0
transform 1 0 12144 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _296_
timestamp 0
transform -1 0 2392 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _297_
timestamp 0
transform 1 0 2944 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 0
transform 1 0 2944 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _299_
timestamp 0
transform 1 0 14904 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _300_
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _301_
timestamp 0
transform 1 0 12604 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 0
transform 1 0 15916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _304_
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _305_
timestamp 0
transform 1 0 4784 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _306_
timestamp 0
transform 1 0 2484 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 0
transform 1 0 2760 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _308_
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _310_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _311_
timestamp 0
transform 1 0 5796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _312_
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _313_
timestamp 0
transform 1 0 10212 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 0
transform 1 0 4416 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _315_
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _316_
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _317_
timestamp 0
transform 1 0 15548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _318_
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _319_
timestamp 0
transform 1 0 7452 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 0
transform 1 0 8648 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _321_
timestamp 0
transform 1 0 12328 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _322_
timestamp 0
transform 1 0 11500 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _323_
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _324_
timestamp 0
transform 1 0 7912 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _325_
timestamp 0
transform 1 0 14444 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _326_
timestamp 0
transform 1 0 5244 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _327_
timestamp 0
transform 1 0 15180 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _328_
timestamp 0
transform 1 0 5244 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _329_
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 0
transform 1 0 9292 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 0
transform 1 0 5520 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _332_
timestamp 0
transform 1 0 10212 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _333_
timestamp 0
transform -1 0 14996 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _334_
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _335_
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _336_
timestamp 0
transform 1 0 2944 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _337_
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _338_
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _339_
timestamp 0
transform 1 0 9660 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _340_
timestamp 0
transform 1 0 14260 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _341_
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _342_
timestamp 0
transform 1 0 4232 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _343_
timestamp 0
transform 1 0 13340 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _344_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _345_
timestamp 0
transform 1 0 12972 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _346_
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_4  _347_
timestamp 0
transform 1 0 2760 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _348_
timestamp 0
transform 1 0 2668 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _349_
timestamp 0
transform 1 0 15364 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _350_
timestamp 0
transform 1 0 14352 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _351_
timestamp 0
transform 1 0 7452 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _352_
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _353_
timestamp 0
transform 1 0 11500 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _354_
timestamp 0
transform 1 0 10764 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _355_
timestamp 0
transform 1 0 2392 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _356_
timestamp 0
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _357_
timestamp 0
transform 1 0 13340 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _358_
timestamp 0
transform 1 0 14812 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _359_
timestamp 0
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _360_
timestamp 0
transform 1 0 7912 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _361_
timestamp 0
transform 1 0 9568 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _362_
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _363_
timestamp 0
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _364_
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _365_
timestamp 0
transform 1 0 11500 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _366_
timestamp 0
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _367_
timestamp 0
transform 1 0 5612 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _368_
timestamp 0
transform 1 0 12604 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _369_
timestamp 0
transform 1 0 10764 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _370_
timestamp 0
transform 1 0 15732 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _371_
timestamp 0
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _372_
timestamp 0
transform 1 0 15824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 0
transform 1 0 5612 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _374_
timestamp 0
transform 1 0 7268 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _376_
timestamp 0
transform 1 0 3772 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _377_
timestamp 0
transform 1 0 5244 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _378_
timestamp 0
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _379_
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 0
transform 1 0 15548 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _381_
timestamp 0
transform 1 0 4600 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _382_
timestamp 0
transform 1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _383_
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _384_
timestamp 0
transform 1 0 14996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _385_
timestamp 0
transform 1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 0
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _387_
timestamp 0
transform 1 0 10120 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _388_
timestamp 0
transform 1 0 9292 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _389_
timestamp 0
transform 1 0 15088 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _390_
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _391_
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _392_
timestamp 0
transform 1 0 2760 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 0
transform 1 0 9016 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _394_
timestamp 0
transform 1 0 10396 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _395_
timestamp 0
transform 1 0 13340 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _396_
timestamp 0
transform 1 0 15088 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _397_
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _398_
timestamp 0
transform 1 0 12604 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _399_
timestamp 0
transform 1 0 10764 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _400_
timestamp 0
transform 1 0 15364 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _401_
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _402_
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _403_
timestamp 0
transform 1 0 6440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _404_
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _405_
timestamp 0
transform 1 0 15640 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _406_
timestamp 0
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _407_
timestamp 0
transform 1 0 1840 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _408_
timestamp 0
transform 1 0 14076 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _409_
timestamp 0
transform 1 0 13984 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _410_
timestamp 0
transform 1 0 4876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _411_
timestamp 0
transform 1 0 2760 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _412_
timestamp 0
transform 1 0 2024 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _414_
timestamp 0
transform 1 0 9844 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _415_
timestamp 0
transform 1 0 7728 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _416_
timestamp 0
transform 1 0 2944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp 0
transform 1 0 13340 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _418_
timestamp 0
transform 1 0 12328 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _419_
timestamp 0
transform 1 0 12696 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _420_
timestamp 0
transform 1 0 14996 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _421_
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _422_
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _423_
timestamp 0
transform 1 0 6624 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _424_
timestamp 0
transform 1 0 3588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _425_
timestamp 0
transform -1 0 15640 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 0
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _427_
timestamp 0
transform 1 0 1564 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _428_
timestamp 0
transform 1 0 2116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _429_
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _430_
timestamp 0
transform 1 0 8188 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _431_
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _432_
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _433_
timestamp 0
transform 1 0 8004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _434_
timestamp 0
transform 1 0 10120 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _435_
timestamp 0
transform 1 0 15088 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _436_
timestamp 0
transform 1 0 13248 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _437_
timestamp 0
transform 1 0 3956 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _438_
timestamp 0
transform 1 0 7912 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _440_
timestamp 0
transform 1 0 11684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _441_
timestamp 0
transform 1 0 9108 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _442_
timestamp 0
transform 1 0 7084 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _443_
timestamp 0
transform 1 0 12512 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _444_
timestamp 0
transform 1 0 10580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _445_
timestamp 0
transform 1 0 15364 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _446_
timestamp 0
transform 1 0 6900 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _447_
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _448_
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _449_
timestamp 0
transform 1 0 9476 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _450_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _451_
timestamp 0
transform 1 0 7452 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _452_
timestamp 0
transform 1 0 9844 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _453_
timestamp 0
transform 1 0 7360 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _454_
timestamp 0
transform 1 0 11408 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _455_
timestamp 0
transform 1 0 13892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _456_
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _457_
timestamp 0
transform 1 0 14996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _458_
timestamp 0
transform 1 0 7820 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _459_
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _460_
timestamp 0
transform 1 0 10396 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _461_
timestamp 0
transform 1 0 15456 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _462_
timestamp 0
transform 1 0 15088 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _463_
timestamp 0
transform 1 0 15180 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _464_
timestamp 0
transform 1 0 15088 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _465_
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _466_
timestamp 0
transform 1 0 12972 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _467_
timestamp 0
transform 1 0 11592 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _468_
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _469_
timestamp 0
transform 1 0 12328 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _470_
timestamp 0
transform 1 0 14904 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _471_
timestamp 0
transform 1 0 14904 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _472_
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _473_
timestamp 0
transform 1 0 12328 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _474_
timestamp 0
transform 1 0 13156 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _475_
timestamp 0
transform 1 0 13800 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _476_
timestamp 0
transform 1 0 12420 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _477_
timestamp 0
transform 1 0 1656 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _478_
timestamp 0
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _479_
timestamp 0
transform 1 0 5152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _480_
timestamp 0
transform 1 0 14352 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _481_
timestamp 0
transform 1 0 1564 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _482_
timestamp 0
transform 1 0 2668 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _483_
timestamp 0
transform 1 0 13524 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _484_
timestamp 0
transform 1 0 6164 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _485_
timestamp 0
transform 1 0 8004 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _486_
timestamp 0
transform 1 0 11592 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _487_
timestamp 0
transform 1 0 15732 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _488_
timestamp 0
transform 1 0 11500 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _489_
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _490_
timestamp 0
transform 1 0 2208 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _491_
timestamp 0
transform 1 0 10764 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _492_
timestamp 0
transform 1 0 6532 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _493_
timestamp 0
transform 1 0 4416 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _495_
timestamp 0
transform 1 0 11500 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _496_
timestamp 0
transform 1 0 4416 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _497_
timestamp 0
transform 1 0 13340 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 0
transform 1 0 6992 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 0
transform 1 0 6072 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _500_
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _501_
timestamp 0
transform 1 0 4232 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 0
transform 1 0 7360 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _505_
timestamp 0
transform 1 0 9200 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _508_
timestamp 0
transform 1 0 11500 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 0
transform 1 0 7084 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _510_
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _511_
timestamp 0
transform 1 0 9660 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _512_
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _513_
timestamp 0
transform 1 0 1472 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _515_
timestamp 0
transform 1 0 1564 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _516_
timestamp 0
transform 1 0 1472 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _517_
timestamp 0
transform 1 0 1840 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp 0
transform 1 0 1472 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _519_
timestamp 0
transform 1 0 3772 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _520_
timestamp 0
transform 1 0 2576 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _521_
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _522_
timestamp 0
transform 1 0 1840 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _523_
timestamp 0
transform 1 0 4232 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _524_
timestamp 0
transform 1 0 1932 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _525_
timestamp 0
transform 1 0 1840 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _526_
timestamp 0
transform 1 0 2576 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _527_
timestamp 0
transform 1 0 1840 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _528_
timestamp 0
transform 1 0 4416 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _529_
timestamp 0
transform 1 0 3772 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _530_
timestamp 0
transform 1 0 1840 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _531_
timestamp 0
transform 1 0 3772 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _532_
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _533_
timestamp 0
transform 1 0 1472 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _534_
timestamp 0
transform 1 0 2576 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _535_
timestamp 0
transform 1 0 1472 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _536_
timestamp 0
transform 1 0 3772 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _537_
timestamp 0
transform 1 0 1472 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _538_
timestamp 0
transform 1 0 4416 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _539_
timestamp 0
transform 1 0 4416 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _540_
timestamp 0
transform 1 0 2576 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _541_
timestamp 0
transform 1 0 2576 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _542_
timestamp 0
transform 1 0 9660 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _543_
timestamp 0
transform 1 0 1472 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _544_
timestamp 0
transform 1 0 4416 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _545_
timestamp 0
transform 1 0 1564 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _546_
timestamp 0
transform 1 0 2024 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _547_
timestamp 0
transform 1 0 1472 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _548_
timestamp 0
transform 1 0 1472 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _549_
timestamp 0
transform 1 0 2208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _550_
timestamp 0
transform 1 0 2944 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _551_
timestamp 0
transform 1 0 3496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _552_
timestamp 0
transform 1 0 2208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _553_
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_0.int_memory_1.GATES_12.result
timestamp 0
transform 1 0 9200 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_0.int_memory_1.GATES_13.result
timestamp 0
transform 1 0 6624 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_0.int_memory_1.GATES_14.result
timestamp 0
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_0.int_memory_1.GATES_15.result
timestamp 0
transform 1 0 8372 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_0.int_memory_1.GATES_16.result
timestamp 0
transform 1 0 8832 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_0.int_memory_1.GATES_17.result
timestamp 0
transform 1 0 9292 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__045_
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__046_
timestamp 0
transform 1 0 9200 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__063_
timestamp 0
transform 1 0 9292 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__220_
timestamp 0
transform 1 0 6992 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__222_
timestamp 0
transform 1 0 8004 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_io_in[0]
timestamp 0
transform 1 0 7912 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_0.int_memory_1.GATES_12.result
timestamp 0
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_0.int_memory_1.GATES_13.result
timestamp 0
transform 1 0 4784 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_0.int_memory_1.GATES_14.result
timestamp 0
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_0.int_memory_1.GATES_15.result
timestamp 0
transform 1 0 4048 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_0.int_memory_1.GATES_16.result
timestamp 0
transform 1 0 5244 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_0.int_memory_1.GATES_17.result
timestamp 0
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__045_
timestamp 0
transform 1 0 10212 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__046_
timestamp 0
transform 1 0 5244 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__063_
timestamp 0
transform 1 0 5244 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__220_
timestamp 0
transform 1 0 5244 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__222_
timestamp 0
transform 1 0 5244 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_io_in[0]
timestamp 0
transform 1 0 4048 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_0.int_memory_1.GATES_12.result
timestamp 0
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_0.int_memory_1.GATES_13.result
timestamp 0
transform 1 0 6624 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_0.int_memory_1.GATES_14.result
timestamp 0
transform 1 0 7820 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_0.int_memory_1.GATES_15.result
timestamp 0
transform 1 0 7820 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_0.int_memory_1.GATES_16.result
timestamp 0
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_0.int_memory_1.GATES_17.result
timestamp 0
transform 1 0 6624 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__045_
timestamp 0
transform 1 0 12788 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__046_
timestamp 0
transform 1 0 10396 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__063_
timestamp 0
transform 1 0 6624 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__220_
timestamp 0
transform 1 0 5244 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__222_
timestamp 0
transform 1 0 9292 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_io_in[0]
timestamp 0
transform 1 0 7820 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform -1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform 1 0 15640 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform 1 0 9016 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 0
transform 1 0 8188 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 0
transform 1 0 14720 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform 1 0 11500 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater8
timestamp 0
transform 1 0 15272 0 -1 16320
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 688 400 808 0 FreeSans 600 0 0 0 io_in[0]
port 1 nsew
flabel metal3 s 0 2184 400 2304 0 FreeSans 600 0 0 0 io_in[1]
port 2 nsew
flabel metal3 s 0 3680 400 3800 0 FreeSans 600 0 0 0 io_in[2]
port 3 nsew
flabel metal3 s 0 5176 400 5296 0 FreeSans 600 0 0 0 io_in[3]
port 4 nsew
flabel metal3 s 0 6672 400 6792 0 FreeSans 600 0 0 0 io_in[4]
port 5 nsew
flabel metal3 s 0 8168 400 8288 0 FreeSans 600 0 0 0 io_in[5]
port 6 nsew
flabel metal3 s 0 9664 400 9784 0 FreeSans 600 0 0 0 io_in[6]
port 7 nsew
flabel metal3 s 0 11160 400 11280 0 FreeSans 600 0 0 0 io_in[7]
port 8 nsew
flabel metal3 s 0 12656 400 12776 0 FreeSans 600 0 0 0 io_out[0]
port 9 nsew
flabel metal3 s 0 14152 400 14272 0 FreeSans 600 0 0 0 io_out[1]
port 10 nsew
flabel metal3 s 0 15648 400 15768 0 FreeSans 600 0 0 0 io_out[2]
port 11 nsew
flabel metal3 s 0 17144 400 17264 0 FreeSans 600 0 0 0 io_out[3]
port 12 nsew
flabel metal3 s 0 18640 400 18760 0 FreeSans 600 0 0 0 io_out[4]
port 13 nsew
flabel metal3 s 0 20136 400 20256 0 FreeSans 600 0 0 0 io_out[5]
port 14 nsew
flabel metal3 s 0 21632 400 21752 0 FreeSans 600 0 0 0 io_out[6]
port 15 nsew
flabel metal3 s 0 23128 400 23248 0 FreeSans 600 0 0 0 io_out[7]
port 16 nsew
flabel metal4 s 2918 1040 3238 22896 0 FreeSans 2400 90 0 0 vccd1
port 17 nsew
flabel metal4 s 6866 1040 7186 22896 0 FreeSans 2400 90 0 0 vccd1
port 17 nsew
flabel metal4 s 10814 1040 11134 22896 0 FreeSans 2400 90 0 0 vccd1
port 17 nsew
flabel metal4 s 14762 1040 15082 22896 0 FreeSans 2400 90 0 0 vccd1
port 17 nsew
flabel metal4 s 4892 1040 5212 22896 0 FreeSans 2400 90 0 0 vssd1
port 18 nsew
flabel metal4 s 8840 1040 9160 22896 0 FreeSans 2400 90 0 0 vssd1
port 18 nsew
flabel metal4 s 12788 1040 13108 22896 0 FreeSans 2400 90 0 0 vssd1
port 18 nsew
<< properties >>
string FIXED_BBOX 0 0 18000 24000
<< end >>
